//: version "1.8.7"

module HA(C, S, B, A);
//: interface  /sz:(148, 128) /bd:[ Li0>B(102/128) Li1>A(35/128) Ro0<C(103/128) Ro1<S(38/128) ]
input B;    //: /sn:0 {0}(197,310)(262,310)(262,284)(288,284){1}
//: {2}(292,284)(337,284){3}
//: {4}(290,286)(290,332)(343,332){5}
input A;    //: /sn:0 {0}(198,279)(304,279){1}
//: {2}(308,279)(337,279){3}
//: {4}(306,281)(306,327)(343,327){5}
output C;    //: /sn:0 /dp:1 {0}(364,330)(448,330){1}
output S;    //: /sn:0 /dp:1 {0}(358,282)(437,282)(437,281)(447,281){1}
//: enddecls

  xor g4 (.I0(A), .I1(B), .Z(S));   //: @(348,282) /sn:0 /delay:" 6" /w:[ 3 3 0 ]
  //: output g3 (C) @(445,330) /sn:0 /w:[ 1 ]
  //: output g2 (S) @(444,281) /sn:0 /w:[ 1 ]
  //: input g1 (B) @(195,310) /sn:0 /w:[ 0 ]
  //: joint g6 (A) @(306, 279) /w:[ 2 -1 1 4 ]
  //: joint g7 (B) @(290, 284) /w:[ 2 -1 1 4 ]
  and g5 (.I0(A), .I1(B), .Z(C));   //: @(354,330) /sn:0 /delay:" 5" /w:[ 5 5 0 ]
  //: input g0 (A) @(196,279) /sn:0 /w:[ 0 ]

endmodule

module main;    //: root_module
wire w4;    //: /sn:0 {0}(654,365)(717,365){1}
wire w0;    //: /sn:0 {0}(449,297)(504,297){1}
wire w1;    //: /sn:0 {0}(449,364)(504,364){1}
wire w5;    //: /sn:0 {0}(654,300)(717,300){1}
//: enddecls

  led g4 (.I(w5));   //: @(724,300) /sn:0 /R:3 /w:[ 1 ] /type:3
  led g3 (.I(w4));   //: @(724,365) /sn:0 /R:3 /w:[ 1 ] /type:3
  HA g2 (.A(w0), .B(w1), .S(w5), .C(w4));   //: @(505, 262) /sz:(148, 128) /sn:0 /p:[ Li0>1 Li1>1 Ro0<0 Ro1<0 ]
  //: switch g1 (w1) @(432,364) /sn:0 /w:[ 0 ] /st:0
  //: switch g0 (w0) @(432,297) /sn:0 /w:[ 0 ] /st:0

endmodule
