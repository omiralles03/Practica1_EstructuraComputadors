//: version "1.8.7"

module FA(Cin, B, S, Cout, A);
//: interface  /sz:(100, 90) /bd:[ Ti0>A(31/100) Ti1>B(74/100) Li0>Cin(43/90) Ri0>S(30/90) Ri1>Cout(69/90) ]
input B;    //: /sn:0 {0}(150,65)(150,107){1}
//: {2}(152,109)(188,109){3}
//: {4}(150,111)(150,159){5}
//: {6}(152,161)(187,161){7}
//: {8}(150,163)(150,182)(187,182){9}
input A;    //: /sn:0 {0}(132,65)(132,102){1}
//: {2}(134,104)(188,104){3}
//: {4}(132,106)(132,128){5}
//: {6}(134,130)(188,130){7}
//: {8}(132,132)(132,156)(187,156){9}
input Cin;    //: /sn:0 {0}(168,65)(168,118){1}
//: {2}(170,120)(259,120)(259,111)(278,111){3}
//: {4}(168,122)(168,133){5}
//: {6}(170,135)(188,135){7}
//: {8}(168,137)(168,187)(187,187){9}
output Cout;    //: /sn:0 /dp:1 {0}(301,149)(340,149){1}
output S;    //: /sn:0 /dp:1 {0}(299,109)(340,109){1}
wire w20;    //: /sn:0 {0}(208,159)(225,159)(225,148)(234,148){1}
wire w8;    //: /sn:0 {0}(208,185)(262,185)(262,151)(280,151){1}
wire w14;    //: /sn:0 {0}(255,146)(280,146){1}
wire w2;    //: /sn:0 {0}(209,106)(278,106){1}
wire w11;    //: /sn:0 {0}(209,133)(225,133)(225,143)(234,143){1}
//: enddecls

  xor g4 (.I0(w2), .I1(Cin), .Z(S));   //: @(289,109) /sn:0 /delay:" 4" /w:[ 1 3 0 ]
  or g8 (.I0(w14), .I1(w8), .Z(Cout));   //: @(291,149) /sn:0 /delay:" 3" /w:[ 1 1 0 ]
  xor g3 (.I0(B), .I1(A), .Z(w2));   //: @(199,106) /sn:0 /delay:" 4" /w:[ 3 3 0 ]
  //: joint g16 (B) @(150, 109) /w:[ 2 1 -1 4 ]
  //: joint g17 (A) @(132, 104) /w:[ 2 1 -1 4 ]
  //: input g2 (Cin) @(168,63) /sn:0 /R:3 /w:[ 0 ]
  //: input g1 (B) @(150,63) /sn:0 /R:3 /w:[ 0 ]
  //: output g10 (S) @(337,109) /sn:0 /w:[ 1 ]
  and g6 (.I0(A), .I1(Cin), .Z(w11));   //: @(199,133) /sn:0 /delay:" 3" /w:[ 7 7 0 ]
  or g7 (.I0(w11), .I1(w20), .Z(w14));   //: @(245,146) /sn:0 /delay:" 3" /w:[ 1 1 0 ]
  and g9 (.I0(A), .I1(B), .Z(w20));   //: @(198,159) /sn:0 /delay:" 3" /w:[ 9 7 0 ]
  //: joint g12 (B) @(150, 161) /w:[ 6 5 -1 8 ]
  and g5 (.I0(B), .I1(Cin), .Z(w8));   //: @(198,185) /sn:0 /delay:" 3" /w:[ 9 9 0 ]
  //: output g11 (Cout) @(337,149) /sn:0 /w:[ 1 ]
  //: joint g14 (A) @(132, 130) /w:[ 6 5 -1 8 ]
  //: input g0 (A) @(132,63) /sn:0 /R:3 /w:[ 0 ]
  //: joint g15 (Cin) @(168, 120) /w:[ 2 1 -1 4 ]
  //: joint g13 (Cin) @(168, 135) /w:[ 6 5 -1 8 ]

endmodule

module main;    //: root_module
wire [3:0] w6;    //: /sn:0 {0}(681,207)(665,207)(665,241){1}
wire w3;    //: /sn:0 {0}(560,281)(594,281){1}
wire w1;    //: /sn:0 {0}(693,283)(722,283){1}
wire [3:0] w2;    //: /sn:0 {0}(644,353)(644,326){1}
wire [3:0] w5;    //: /sn:0 {0}(608,207)(624,207)(624,241){1}
//: enddecls

  //: switch g4 (w3) @(543,281) /sn:0 /w:[ 0 ] /st:1
  led g3 (.I(w2));   //: @(644,360) /sn:0 /R:2 /w:[ 0 ] /type:2
  //: dip g2 (w6) @(719,207) /sn:0 /R:3 /w:[ 0 ] /st:3
  //: dip g1 (w5) @(570,207) /sn:0 /R:1 /w:[ 0 ] /st:11
  led g5 (.I(w1));   //: @(729,283) /sn:0 /R:3 /w:[ 1 ] /type:2
  CPA_4b g0 (.B(w6), .A(w5), .Cin(w3), .S(w2), .Cout(w1));   //: @(595, 242) /sz:(97, 83) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>1 Bo0<1 Ro0<0 ]

endmodule

module CPA_4b(S, Cin, Cout, B, A);
//: interface  /sz:(97, 83) /bd:[ Ti0>A[3:0](29/97) Ti1>B[3:0](70/97) Li0>Cin(39/83) Bo0<S[3:0](49/97) Ro0<Cout(41/83) ]
input [3:0] B;    //: /sn:0 {0}(298,170)(413,170){1}
//: {2}(414,170)(550,170){3}
//: {4}(551,170)(679,170){5}
//: {6}(680,170)(816,170){7}
//: {8}(817,170)(900,170){9}
input [3:0] A;    //: /sn:0 {0}(896,147)(774,147){1}
//: {2}(773,147)(637,147){3}
//: {4}(636,147)(508,147){5}
//: {6}(507,147)(371,147){7}
//: {8}(370,147)(299,147){9}
input Cin;    //: /sn:0 {0}(295,231)(343,231){1}
output Cout;    //: /sn:0 /dp:1 {0}(848,235)(911,235){1}
output [3:0] S;    //: /sn:0 {0}(877,326)(922,326){1}
wire w13;    //: /sn:0 {0}(637,201)(637,151){1}
wire w16;    //: /sn:0 {0}(658,292)(658,321)(871,321){1}
wire w7;    //: /sn:0 {0}(817,202)(817,174){1}
wire w4;    //: /sn:0 {0}(371,199)(371,151){1}
wire w0;    //: /sn:0 {0}(551,200)(551,174){1}
wire w3;    //: /sn:0 /dp:1 {0}(871,331)(529,331)(529,291){1}
wire w10;    //: /sn:0 {0}(680,201)(680,174){1}
wire w1;    //: /sn:0 {0}(508,200)(508,151){1}
wire w8;    //: /sn:0 /dp:1 {0}(480,232)(445,232){1}
wire w14;    //: /sn:0 /dp:1 {0}(609,233)(582,233){1}
wire w2;    //: /sn:0 {0}(414,199)(414,174){1}
wire w11;    //: /sn:0 /dp:1 {0}(392,290)(392,341)(871,341){1}
wire w15;    //: /sn:0 /dp:1 {0}(746,234)(711,234){1}
wire w5;    //: /sn:0 /dp:1 {0}(871,311)(795,311)(795,293){1}
wire w9;    //: /sn:0 {0}(774,202)(774,151){1}
//: enddecls

  //: output g8 (S) @(919,326) /sn:0 /w:[ 1 ]
  FA g4 (.A(w4), .B(w2), .Cin(Cin), .S(w11), .Cout(w8));   //: @(344, 200) /sz:(100, 89) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>1 Bo0<0 Ro0<1 ]
  tran g16(.Z(w9), .I(A[3]));   //: @(774,145) /sn:0 /R:1 /w:[ 1 2 1 ] /ss:1
  //: input g3 (Cin) @(293,231) /sn:0 /w:[ 0 ]
  tran g17(.Z(w7), .I(B[3]));   //: @(817,168) /sn:0 /R:1 /w:[ 1 7 8 ] /ss:1
  //: output g2 (Cout) @(908,235) /sn:0 /w:[ 1 ]
  //: input g1 (B) @(296,170) /sn:0 /w:[ 0 ]
  tran g10(.Z(w4), .I(A[0]));   //: @(371,145) /sn:0 /R:1 /w:[ 1 8 7 ] /ss:1
  FA g6 (.A(w13), .B(w10), .Cin(w14), .S(w16), .Cout(w15));   //: @(610, 202) /sz:(100, 89) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>0 Bo0<0 Ro0<1 ]
  concat g9 (.I0(w11), .I1(w3), .I2(w16), .I3(w5), .Z(S));   //: @(876,326) /sn:0 /w:[ 1 0 1 0 0 ] /dr:0
  FA g7 (.A(w9), .B(w7), .Cin(w15), .S(w5), .Cout(Cout));   //: @(747, 203) /sz:(100, 89) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>0 Bo0<1 Ro0<0 ]
  tran g12(.Z(w1), .I(A[1]));   //: @(508,145) /sn:0 /R:1 /w:[ 1 6 5 ] /ss:1
  tran g14(.Z(w13), .I(A[2]));   //: @(637,145) /sn:0 /R:1 /w:[ 1 4 3 ] /ss:1
  tran g11(.Z(w2), .I(B[0]));   //: @(414,168) /sn:0 /R:1 /w:[ 1 1 2 ] /ss:1
  FA g5 (.A(w1), .B(w0), .Cin(w8), .S(w3), .Cout(w14));   //: @(481, 201) /sz:(100, 89) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>0 Bo0<1 Ro0<1 ]
  tran g15(.Z(w10), .I(B[2]));   //: @(680,168) /sn:0 /R:1 /w:[ 1 5 6 ] /ss:1
  //: input g0 (A) @(297,147) /sn:0 /w:[ 9 ]
  tran g13(.Z(w0), .I(B[1]));   //: @(551,168) /sn:0 /R:1 /w:[ 1 3 4 ] /ss:1

endmodule
