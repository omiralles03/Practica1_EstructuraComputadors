//: version "1.8.7"

module RPA4(B, S, A);
//: interface  /sz:(119, 111) /bd:[ Ti0>A[3:0](22/119) Ti1>B[3:0](105/119) Bo0<S[7:0](58/119) ]
input [3:0] B;    //: /sn:0 /dp:1 {0}(155,208)(123,208){1}
input [3:0] A;    //: /sn:0 /dp:11 {0}(413,279)(444,279){1}
//: {2}(445,279)(538,279)(538,277)(646,277){3}
//: {4}(647,277)(709,277)(709,278)(755,278){5}
//: {6}(756,278)(788,278)(788,276)(808,276){7}
//: {8}(809,276)(1056,276)(1056,343)(1267,343){9}
//: {10}(1271,343)(1433,343)(1433,342)(1443,342){11}
//: {12}(1269,341)(1269,54)(687,54){13}
//: {14}(686,54)(651,54)(651,53)(628,53){15}
//: {16}(627,53)(578,53){17}
//: {18}(577,53)(499,53){19}
//: {20}(498,53)(454,53){21}
//: {22}(453,53)(404,53)(404,54)(299,54){23}
//: {24}(298,54)(275,54){25}
//: {26}(274,54)(229,54){27}
//: {28}(228,54)(193,54){29}
//: {30}(1269,345)(1269,467)(1073,467){31}
//: {32}(1072,467)(914,467){33}
//: {34}(913,467)(903,467)(903,465)(793,465){35}
//: {36}(792,465)(725,465)(725,464)(564,464){37}
//: {38}(563,464)(539,464){39}
output [7:0] S;    //: /sn:0 /dp:1 {0}(1324,723)(1391,723)(1391,724)(1397,724){1}
wire w13;    //: /sn:0 {0}(301,153)(301,215)(308,215){1}
wire w16;    //: /sn:0 {0}(445,283)(445,342){1}
wire w6;    //: /sn:0 {0}(687,58)(687,82)(682,82)(682,138){1}
wire w58;    //: /sn:0 {0}(1075,549)(1075,571){1}
wire w7;    //: /sn:0 {0}(578,57)(578,86){1}
wire w65;    //: /sn:0 /dp:1 {0}(1318,738)(897,738)(897,656){1}
wire w50;    //: /sn:0 {0}(1077,528)(1077,503)(937,503){1}
//: {2}(933,503)(923,503)(923,504)(812,504){3}
//: {4}(808,504)(696,504)(696,505)(579,505){5}
//: {6}(575,505)(181,505)(181,223)(161,223){7}
//: {8}(577,507)(577,514)(570,514)(570,524){9}
//: {10}(810,506)(810,531)(798,531)(798,541){11}
//: {12}(935,505)(935,531)(926,531)(926,539){13}
wire w34;    //: /sn:0 {0}(809,280)(809,297)(857,297)(857,322){1}
wire w59;    //: /sn:0 /dp:1 {0}(1318,708)(554,708)(554,410)(542,410){1}
wire w25;    //: /sn:0 {0}(774,233)(914,233)(914,352)(807,352)(807,367){1}
wire w4;    //: /sn:0 {0}(454,57)(454,83){1}
wire w62;    //: /sn:0 /dp:1 {0}(1318,718)(726,718)(726,587)(680,587){1}
wire w56;    //: /sn:0 {0}(815,628)(849,628)(849,627)(858,627){1}
wire w22;    //: /sn:0 {0}(517,229)(570,229){1}
wire w36;    //: /sn:0 {0}(667,405)(689,405)(689,404)(701,404){1}
wire w0;    //: /sn:0 {0}(161,193)(180,193)(180,74)(234,74){1}
//: {2}(238,74)(256,74)(256,72)(266,72){3}
//: {4}(270,72)(385,72)(385,71)(456,71){5}
//: {6}(460,71)(569,71)(569,72)(581,72){7}
//: {8}(585,72)(732,72){9}
//: {10}(583,74)(583,86){11}
//: {12}(458,73)(458,78)(459,78)(459,83){13}
//: {14}(268,74)(268,97)(270,97)(270,98){15}
//: {16}(236,76)(236,381)(234,381)(234,395){17}
wire w20;    //: /sn:0 {0}(392,225)(411,225)(411,227)(431,227){1}
wire w29;    //: /sn:0 {0}(581,107)(581,174)(580,174)(580,185){1}
wire w42;    //: /sn:0 {0}(862,322)(862,306)(769,306){1}
//: {2}(765,306)(653,306){3}
//: {4}(649,306)(533,306)(533,318)(452,318){5}
//: {6}(448,318)(200,318)(200,213)(161,213){7}
//: {8}(450,320)(450,342){9}
//: {10}(651,308)(651,321){11}
//: {12}(767,308)(767,312)(761,312)(761,326){13}
wire w37;    //: /sn:0 {0}(649,342)(649,353){1}
wire w12;    //: /sn:0 {0}(272,119)(272,187)(308,187){1}
wire w18;    //: /sn:0 {0}(651,235)(689,235)(689,224)(699,224){1}
wire w10;    //: /sn:0 {0}(231,416)(231,688)(1318,688){1}
wire w23;    //: /sn:0 {0}(628,57)(628,96)(626,96)(626,134){1}
wire w63;    //: /sn:0 {0}(796,562)(796,569)(798,569)(798,577){1}
wire w54;    //: /sn:0 {0}(564,468)(564,498)(565,498)(565,524){1}
wire w24;    //: /sn:0 {0}(774,199)(863,199)(863,258)(722,258)(722,363){1}
wire w21;    //: /sn:0 {0}(471,258)(471,312)(461,312)(461,367)(471,367){1}
wire w1;    //: /sn:0 {0}(161,203)(205,203)(205,115)(302,115){1}
//: {2}(306,115)(404,115)(404,116)(502,116){3}
//: {4}(506,116)(629,116){5}
//: {6}(633,116)(641,116)(641,117)(691,117){7}
//: {8}(695,117)(780,117){9}
//: {10}(693,119)(693,129)(687,129)(687,138){11}
//: {12}(631,118)(631,134){13}
//: {14}(504,118)(504,127)(503,127)(503,129){15}
//: {16}(304,117)(304,132){17}
wire w31;    //: /sn:0 {0}(542,395)(551,395)(551,399)(581,399){1}
wire w32;    //: /sn:0 {0}(756,282)(756,326){1}
wire w68;    //: /sn:0 {0}(746,577)(746,489)(736,489)(736,430){1}
wire w53;    //: /sn:0 {0}(1092,619)(1212,619)(1212,758)(1318,758){1}
wire w8;    //: /sn:0 {0}(275,58)(275,98){1}
wire w52;    //: /sn:0 {0}(914,471)(914,536)(921,536)(921,539){1}
wire w27;    //: /sn:0 {0}(629,155)(629,166)(634,166)(634,185){1}
wire w44;    //: /sn:0 {0}(874,410)(1047,410)(1047,450)(1021,450)(1021,571){1}
wire w17;    //: /sn:0 {0}(609,257)(609,287)(592,287)(592,353){1}
wire w33;    //: /sn:0 {0}(448,363)(448,407)(471,407){1}
wire w35;    //: /sn:0 {0}(621,434)(621,558)(574,558)(574,585)(595,585){1}
wire w28;    //: /sn:0 {0}(685,159)(685,197)(699,197){1}
wire w49;    //: /sn:0 {0}(1073,471)(1073,499)(1072,499)(1072,528){1}
wire w14;    //: /sn:0 {0}(500,150)(500,163)(499,163)(499,176){1}
wire w45;    //: /sn:0 {0}(860,343)(860,350)(858,350)(858,367){1}
wire w11;    //: /sn:0 {0}(299,58)(299,132){1}
wire w2;    //: /sn:0 {0}(793,469)(793,541){1}
wire w41;    //: /sn:0 {0}(759,347)(759,357)(760,357)(760,363){1}
wire w48;    //: /sn:0 {0}(1318,698)(420,698)(420,189)(392,189){1}
wire w47;    //: /sn:0 {0}(680,628)(726,628)(726,626)(736,626){1}
wire w15;    //: /sn:0 {0}(457,104)(457,134)(442,134)(442,176){1}
wire w5;    //: /sn:0 {0}(499,57)(499,64)(498,64)(498,129){1}
wire w38;    //: /sn:0 {0}(595,621)(567,621)(567,545){1}
wire w61;    //: /sn:0 {0}(941,629)(967,629)(967,617)(1011,617){1}
wire w43;    //: /sn:0 {0}(833,434)(833,550)(869,550)(869,581){1}
wire w64;    //: /sn:0 /dp:1 {0}(1318,728)(773,728)(773,656){1}
wire w26;    //: /sn:0 {0}(647,281)(647,298)(646,298)(646,321){1}
wire w9;    //: /sn:0 {0}(229,58)(229,395){1}
wire w57;    //: /sn:0 {0}(924,560)(924,572)(923,572)(923,581){1}
wire w40;    //: /sn:0 {0}(776,406)(794,406)(794,408)(797,408){1}
wire w51;    //: /sn:0 {0}(1049,646)(1049,748)(1318,748){1}
//: enddecls

  and g44 (.I0(w34), .I1(w42), .Z(w45));   //: @(860,333) /sn:0 /R:3 /delay:" 5" /w:[ 1 0 0 ]
  tran g8(.Z(w8), .I(A[1]));   //: @(275,52) /sn:0 /R:1 /w:[ 0 26 25 ] /ss:1
  tran g4(.Z(w9), .I(A[0]));   //: @(229,52) /sn:0 /R:1 /w:[ 0 28 27 ] /ss:1
  HalfAdder g47 (.b(w38), .a(w35), .c(w47), .s(w62));   //: @(596, 568) /sz:(83, 76) /sn:0 /p:[ Li0>0 Li1>1 Ro0<0 Ro1<1 ]
  //: joint g16 (w0) @(458, 71) /w:[ 6 -1 5 12 ]
  and g3 (.I0(w0), .I1(w9), .Z(w10));   //: @(231,406) /sn:0 /R:3 /delay:" 5" /w:[ 17 1 0 ]
  HalfAdder g26 (.b(w13), .a(w12), .c(w20), .s(w48));   //: @(309, 173) /sz:(82, 66) /sn:0 /p:[ Li0>1 Li1>1 Ro0<0 Ro1<1 ]
  FullAdder g17 (.b(w27), .a(w29), .Cin(w22), .s(w17), .Cout(w18));   //: @(571, 186) /sz:(79, 70) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>1 Bo0<0 Ro0<0 ]
  concat g2 (.I0(w0), .I1(w1), .I2(w42), .I3(w50), .Z(B));   //: @(156,208) /sn:0 /R:2 /w:[ 0 0 7 7 0 ] /dr:0
  tran g30(.Z(w6), .I(A[3]));   //: @(687,52) /sn:0 /R:1 /w:[ 0 14 13 ] /ss:1
  //: joint g23 (w0) @(583, 72) /w:[ 8 -1 7 10 ]
  //: joint g24 (w1) @(631, 116) /w:[ 6 -1 5 12 ]
  FullAdder g39 (.b(w41), .a(w24), .Cin(w36), .s(w68), .Cout(w40));   //: @(702, 364) /sz:(73, 65) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>1 Bo0<1 Ro0<0 ]
  //: input g1 (B) @(121,208) /sn:0 /w:[ 1 ]
  tran g60(.Z(w52), .I(A[2]));   //: @(914,465) /sn:0 /R:1 /w:[ 0 34 33 ] /ss:1
  //: joint g29 (w1) @(693, 117) /w:[ 8 -1 7 10 ]
  and g51 (.I0(w50), .I1(w54), .Z(w38));   //: @(567,535) /sn:0 /R:3 /delay:" 5" /w:[ 9 1 1 ]
  tran g18(.Z(w5), .I(A[1]));   //: @(499,51) /sn:0 /R:1 /w:[ 0 20 19 ] /ss:1
  tran g25(.Z(w23), .I(A[2]));   //: @(628,51) /sn:0 /R:1 /w:[ 0 16 15 ] /ss:1
  tran g10(.Z(w11), .I(A[0]));   //: @(299,52) /sn:0 /R:1 /w:[ 0 24 23 ] /ss:1
  concat g64 (.I0(w10), .I1(w48), .I2(w59), .I3(w62), .I4(w64), .I5(w65), .I6(w51), .I7(w53), .Z(S));   //: @(1323,723) /sn:0 /w:[ 1 0 0 0 0 0 1 1 0 ] /dr:1
  FullAdder g49 (.b(w63), .a(w68), .Cin(w47), .s(w64), .Cout(w56));   //: @(737, 578) /sz:(77, 77) /sn:0 /p:[ Ti0>1 Ti1>0 Li0>1 Bo0<1 Ro0<0 ]
  and g6 (.I0(w8), .I1(w0), .Z(w12));   //: @(272,109) /sn:0 /R:3 /delay:" 5" /w:[ 1 15 0 ]
  FullAdder g50 (.b(w57), .a(w43), .Cin(w56), .s(w65), .Cout(w61));   //: @(859, 582) /sz:(81, 73) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>1 Bo0<1 Ro0<0 ]
  FullAdder g35 (.b(w37), .a(w17), .Cin(w31), .s(w35), .Cout(w36));   //: @(582, 354) /sz:(84, 79) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>1 Bo0<0 Ro0<0 ]
  tran g56(.Z(w2), .I(A[1]));   //: @(793,463) /sn:0 /R:1 /w:[ 0 36 35 ] /ss:1
  and g9 (.I0(w1), .I1(w11), .Z(w13));   //: @(301,143) /sn:0 /R:3 /delay:" 5" /w:[ 17 1 0 ]
  //: joint g7 (w0) @(268, 72) /w:[ 4 -1 3 14 ]
  and g58 (.I0(w52), .I1(w50), .Z(w57));   //: @(924,550) /sn:0 /R:3 /delay:" 5" /w:[ 1 13 0 ]
  tran g22(.Z(w7), .I(A[3]));   //: @(578,51) /sn:0 /R:1 /w:[ 0 18 17 ] /ss:1
  HalfAdder g31 (.b(w33), .a(w21), .c(w31), .s(w59));   //: @(472, 352) /sz:(69, 69) /sn:0 /p:[ Li0>1 Li1>1 Ro0<0 Ro1<1 ]
  //: joint g59 (w50) @(935, 503) /w:[ 1 -1 2 12 ]
  //: joint g33 (w42) @(450, 318) /w:[ 5 -1 6 8 ]
  tran g45(.Z(w34), .I(A[3]));   //: @(809,274) /sn:0 /R:1 /w:[ 0 7 8 ] /ss:1
  and g54 (.I0(w2), .I1(w50), .Z(w63));   //: @(796,552) /sn:0 /R:3 /delay:" 5" /w:[ 1 11 0 ]
  //: joint g41 (w42) @(767, 306) /w:[ 1 -1 2 12 ]
  and g36 (.I0(w26), .I1(w42), .Z(w37));   //: @(649,332) /sn:0 /R:3 /delay:" 5" /w:[ 1 11 0 ]
  and g40 (.I0(w32), .I1(w42), .Z(w41));   //: @(759,337) /sn:0 /R:3 /delay:" 5" /w:[ 1 13 0 ]
  tran g42(.Z(w32), .I(A[2]));   //: @(756,276) /sn:0 /R:1 /w:[ 0 5 6 ] /ss:1
  tran g52(.Z(w54), .I(A[0]));   //: @(564,462) /sn:0 /R:1 /w:[ 0 38 37 ] /ss:1
  and g12 (.I0(w1), .I1(w5), .Z(w14));   //: @(500,140) /sn:0 /R:3 /delay:" 5" /w:[ 15 1 0 ]
  and g28 (.I0(w6), .I1(w1), .Z(w28));   //: @(685,149) /sn:0 /R:3 /delay:" 5" /w:[ 1 11 0 ]
  tran g34(.Z(w16), .I(A[0]));   //: @(445,277) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:1
  //: joint g46 (A) @(1269, 343) /w:[ 10 12 9 30 ]
  and g14 (.I0(w4), .I1(w0), .Z(w15));   //: @(457,94) /sn:0 /R:3 /delay:" 5" /w:[ 1 13 0 ]
  //: joint g5 (w0) @(236, 74) /w:[ 2 -1 1 16 ]
  //: joint g11 (w1) @(304, 115) /w:[ 2 -1 1 16 ]
  and g21 (.I0(w7), .I1(w0), .Z(w29));   //: @(581,97) /sn:0 /R:3 /delay:" 5" /w:[ 1 11 0 ]
  HalfAdder g19 (.b(w18), .a(w28), .c(w25), .s(w24));   //: @(700, 184) /sz:(73, 62) /sn:0 /p:[ Li0>1 Li1>1 Ro0<0 Ro1<0 ]
  and g61 (.I0(w49), .I1(w50), .Z(w58));   //: @(1075,539) /sn:0 /R:3 /delay:" 5" /w:[ 1 0 0 ]
  and g20 (.I0(w23), .I1(w1), .Z(w27));   //: @(629,145) /sn:0 /R:3 /delay:" 5" /w:[ 1 13 0 ]
  and g32 (.I0(w16), .I1(w42), .Z(w33));   //: @(448,353) /sn:0 /R:3 /delay:" 5" /w:[ 1 9 0 ]
  //: output g63 (S) @(1394,724) /sn:0 /w:[ 1 ]
  //: input g0 (A) @(1445,342) /sn:0 /R:2 /w:[ 11 ]
  FullAdder g43 (.b(w45), .a(w25), .Cin(w40), .s(w43), .Cout(w44));   //: @(798, 368) /sz:(75, 65) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>1 Bo0<0 Ro0<0 ]
  tran g15(.Z(w4), .I(A[2]));   //: @(454,51) /sn:0 /R:1 /w:[ 0 22 21 ] /ss:1
  tran g38(.Z(w26), .I(A[1]));   //: @(647,275) /sn:0 /R:1 /w:[ 0 3 4 ] /ss:1
  FullAdder g48 (.a(w44), .b(w58), .Cin(w61), .s(w51), .Cout(w53));   //: @(1012, 572) /sz:(79, 73) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>1 Bo0<0 Ro0<0 ]
  FullAdder g27 (.b(w14), .a(w15), .Cin(w20), .s(w21), .Cout(w22));   //: @(432, 177) /sz:(84, 80) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>1 Bo0<0 Ro0<0 ]
  tran g62(.Z(w49), .I(A[3]));   //: @(1073,465) /sn:0 /R:1 /w:[ 0 32 31 ] /ss:1
  //: joint g37 (w42) @(651, 306) /w:[ 3 -1 4 10 ]
  //: joint g55 (w50) @(810, 504) /w:[ 3 -1 4 10 ]
  //: joint g53 (w50) @(577, 505) /w:[ 5 -1 6 8 ]
  //: joint g13 (w1) @(504, 116) /w:[ 4 -1 3 14 ]

endmodule

module FullAdder(Cin, b, a, s, Cout);
//: interface  /sz:(89, 89) /bd:[ Ti0>a(13/89) Ti1>b(73/89) Li0>Cin(57/89) Bo0<s(44/89) Ro0<Cout(58/89) ]
input b;    //: /sn:0 {0}(172,118)(285,118){1}
input Cin;    //: /sn:0 /dp:1 {0}(450,127)(434,127)(434,208)(453,208){1}
output Cout;    //: /sn:0 /dp:1 {0}(613,235)(677,235){1}
output s;    //: /sn:0 /dp:1 {0}(531,94)(685,94){1}
input a;    //: /sn:0 {0}(171,89)(285,89){1}
wire w3;    //: /sn:0 /dp:1 {0}(592,232)(568,232)(568,129)(531,129){1}
wire w1;    //: /sn:0 {0}(450,92)(366,92){1}
wire w2;    //: /sn:0 {0}(366,127)(412,127)(412,237)(592,237){1}
//: enddecls

  //: input g4 (Cin) @(455,208) /sn:0 /R:2 /w:[ 1 ]
  //: input g3 (b) @(170,118) /sn:0 /w:[ 0 ]
  //: input g2 (a) @(169,89) /sn:0 /w:[ 0 ]
  HalfAdder g1 (.a(w1), .b(Cin), .s(s), .c(w3));   //: @(451, 76) /sz:(79, 66) /sn:0 /p:[ Li0>0 Li1>0 Ro0<0 Ro1<1 ]
  //: output g12 (s) @(682,94) /sn:0 /w:[ 1 ]
  or g5 (.I0(w3), .I1(w2), .Z(Cout));   //: @(603,235) /sn:0 /delay:" 5" /w:[ 0 1 0 ]
  HalfAdder g0 (.a(a), .b(b), .s(w1), .c(w2));   //: @(286, 74) /sz:(79, 66) /sn:0 /p:[ Li0>1 Li1>1 Ro0<1 Ro1<0 ]
  //: output g13 (Cout) @(674,235) /sn:0 /w:[ 1 ]

endmodule

module main;    //: root_module
wire [3:0] B;    //: /sn:0 /dp:1 {0}(604,114)(604,207)(561,207)(561,252){1}
wire [3:0] A;    //: /sn:0 {0}(410,112)(410,205)(478,205)(478,252){1}
wire [7:0] S;    //: /sn:0 {0}(514,365)(514,444){1}
//: enddecls

  led g3 (.I(S));   //: @(514,451) /sn:0 /R:2 /w:[ 1 ] /type:3
  //: dip g2 (B) @(604,104) /sn:0 /w:[ 0 ] /st:5
  //: dip g1 (A) @(410,102) /sn:0 /w:[ 0 ] /st:3
  RPA4 g0 (.B(B), .A(A), .S(S));   //: @(456, 253) /sz:(119, 111) /sn:0 /p:[ Ti0>1 Ti1>1 Bo0<0 ]

endmodule

module HalfAdder(s, b, a, c);
//: interface  /sz:(79, 66) /bd:[ Li0>a(16/66) Li1>b(44/66) Ro0<s(18/66) Ro1<c(53/66) ]
input b;    //: /sn:0 /dp:1 {0}(424,277)(354,277){1}
//: {2}(352,275)(352,226)(426,226){3}
//: {4}(350,277)(302,277){5}
output s;    //: /sn:0 {0}(491,224)(447,224){1}
input a;    //: /sn:0 {0}(301,217)(389,217){1}
//: {2}(393,217)(409,217)(409,221)(426,221){3}
//: {4}(391,219)(391,272)(424,272){5}
output c;    //: /sn:0 /dp:1 {0}(445,275)(495,275){1}
//: enddecls

  //: output g4 (s) @(488,224) /sn:0 /w:[ 0 ]
  //: input g3 (b) @(300,277) /sn:0 /w:[ 5 ]
  //: input g2 (a) @(299,217) /sn:0 /w:[ 0 ]
  and g1 (.I0(a), .I1(b), .Z(c));   //: @(435,275) /sn:0 /delay:" 5" /w:[ 5 0 0 ]
  //: joint g6 (a) @(391, 217) /w:[ 2 -1 1 4 ]
  //: joint g7 (b) @(352, 277) /w:[ 1 2 4 -1 ]
  //: output g5 (c) @(492,275) /sn:0 /w:[ 1 ]
  xor g0 (.I0(a), .I1(b), .Z(s));   //: @(437,224) /sn:0 /delay:" 6" /w:[ 3 3 1 ]

endmodule
