//: version "1.8.7"

module CSA_16b(A, S, Cin, Co, B);
//: interface  /sz:(226, 126) /bd:[ Ti0>B[15:0](136/226) Ti1>A[15:0](58/226) Ri0>Cin(60/126) Lo0<Co(63/126) Bo0<S[15:0](102/226) ]
input [15:0] B;    //: /sn:0 {0}(118,-1)(304,-1){1}
//: {2}(305,-1)(564,-1){3}
//: {4}(565,-1)(837,-1){5}
//: {6}(838,-1)(1104,-1){7}
//: {8}(1105,-1)(1121,-1){9}
input [15:0] A;    //: /sn:0 {0}(1121,-49)(1022,-49){1}
//: {2}(1021,-49)(771,-49){3}
//: {4}(770,-49)(498,-49){5}
//: {6}(497,-49)(248,-49){7}
//: {8}(247,-49)(118,-49){9}
input Cin;    //: /sn:0 {0}(1333,221)(1232,221)(1232,196)(1156,196){1}
output Co;    //: /sn:0 /dp:1 {0}(203,203)(104,203)(104,206)(94,206){1}
output [15:0] S;    //: /sn:0 /dp:1 {0}(37,433)(135,433)(135,445)(145,445){1}
wire w13;    //: /sn:0 {0}(729,203)(620,203)(620,210)(610,210){1}
wire [3:0] w6;    //: /sn:0 /dp:1 {0}(498,-45)(498,127)(497,127)(497,137){1}
wire [3:0] w16;    //: /sn:0 /dp:1 {0}(1105,3)(1105,135)(1106,135)(1106,145){1}
wire [3:0] w3;    //: /sn:0 {0}(1061,284)(1061,430)(151,430){1}
wire [3:0] w0;    //: /sn:0 {0}(774,131)(774,103)(771,103)(771,-45){1}
wire [3:0] w20;    //: /sn:0 {0}(307,131)(307,11)(305,11)(305,3){1}
wire [3:0] w19;    //: /sn:0 {0}(528,281)(528,450)(151,450){1}
wire w18;    //: /sn:0 {0}(452,209)(371,209)(371,204)(361,204){1}
wire [3:0] w24;    //: /sn:0 {0}(279,275)(279,460)(151,460){1}
wire [3:0] w21;    //: /sn:0 {0}(248,131)(248,-45){1}
wire w8;    //: /sn:0 {0}(972,250)(897,250)(897,204)(887,204){1}
wire [3:0] w14;    //: /sn:0 {0}(805,275)(805,500)(441,500)(441,440)(151,440){1}
wire [3:0] w2;    //: /sn:0 /dp:1 {0}(833,131)(833,90)(838,90)(838,3){1}
wire [3:0] w15;    //: /sn:0 /dp:1 {0}(1022,-45)(1022,135)(1026,135)(1026,145){1}
wire [3:0] w5;    //: /sn:0 {0}(565,3)(565,127)(556,127)(556,137){1}
//: enddecls

  //: input g4 (A) @(116,-49) /sn:0 /w:[ 9 ]
  tran g8(.Z(w16), .I(B[3:0]));   //: @(1105,-3) /sn:0 /R:1 /w:[ 0 7 8 ] /ss:1
  tran g16(.Z(w20), .I(B[15:12]));   //: @(305,-3) /sn:0 /R:1 /w:[ 1 1 2 ] /ss:1
  CSA_4bit g3 (.A(w6), .B(w5), .Ci(w13), .Co(w18), .S(w19));   //: @(453, 138) /sz:(156, 142) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  //: output g17 (S) @(40,433) /sn:0 /R:2 /w:[ 0 ]
  CSA_4bit g2 (.A(w0), .B(w2), .Ci(w8), .Co(w13), .S(w14));   //: @(730, 132) /sz:(156, 142) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Lo0<0 Bo0<0 ]
  concat g1 (.I0(w3), .I1(w14), .I2(w19), .I3(w24), .Z(S));   //: @(146,445) /sn:0 /R:2 /w:[ 1 1 1 1 1 ] /dr:0
  tran g10(.Z(w0), .I(A[7:4]));   //: @(771,-51) /sn:0 /R:1 /w:[ 1 4 3 ] /ss:1
  tran g6(.Z(w6), .I(A[11:8]));   //: @(498,-51) /sn:0 /R:1 /w:[ 0 6 5 ] /ss:1
  tran g7(.Z(w15), .I(A[3:0]));   //: @(1022,-51) /sn:0 /R:1 /w:[ 0 2 1 ] /ss:1
  tran g9(.Z(w2), .I(B[7:4]));   //: @(838,-3) /sn:0 /R:1 /w:[ 1 5 6 ] /ss:1
  //: input g12 (Cin) @(1335,221) /sn:0 /R:2 /w:[ 0 ]
  //: output g14 (Co) @(97,206) /sn:0 /R:2 /w:[ 1 ]
  //: input g5 (B) @(116,-1) /sn:0 /w:[ 0 ]
  tran g11(.Z(w5), .I(B[11:8]));   //: @(565,-3) /sn:0 /R:1 /w:[ 0 3 4 ] /ss:1
  tran g15(.Z(w21), .I(A[15:12]));   //: @(248,-51) /sn:0 /R:1 /w:[ 1 8 7 ] /ss:1
  CPA g0 (.B(w16), .A(w15), .Ci(Cin), .Co(w8), .S(w3));   //: @(973, 146) /sz:(182, 137) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  CSA_4bit g13 (.A(w21), .B(w20), .Ci(w18), .Co(Co), .S(w24));   //: @(204, 132) /sz:(156, 142) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Lo0<0 Bo0<0 ]

endmodule

module HA(C, S, B, A);
//: interface  /sz:(148, 128) /bd:[ Li0>A(35/128) Li1>B(102/128) Ro0<S(38/128) Ro1<C(103/128) ]
input B;    //: /sn:0 {0}(197,310)(262,310)(262,284)(288,284){1}
//: {2}(292,284)(337,284){3}
//: {4}(290,286)(290,332)(343,332){5}
input A;    //: /sn:0 {0}(198,279)(304,279){1}
//: {2}(308,279)(337,279){3}
//: {4}(306,281)(306,327)(343,327){5}
output C;    //: /sn:0 /dp:1 {0}(364,330)(448,330){1}
output S;    //: /sn:0 /dp:1 {0}(358,282)(437,282)(437,281)(447,281){1}
//: enddecls

  xor g4 (.I0(A), .I1(B), .Z(S));   //: @(348,282) /sn:0 /delay:" 6" /w:[ 3 3 0 ]
  //: output g3 (C) @(445,330) /sn:0 /w:[ 1 ]
  //: output g2 (S) @(444,281) /sn:0 /w:[ 1 ]
  //: input g1 (B) @(195,310) /sn:0 /w:[ 0 ]
  //: joint g6 (A) @(306, 279) /w:[ 2 -1 1 4 ]
  //: joint g7 (B) @(290, 284) /w:[ 2 -1 1 4 ]
  and g5 (.I0(A), .I1(B), .Z(C));   //: @(354,330) /sn:0 /delay:" 5" /w:[ 5 5 0 ]
  //: input g0 (A) @(196,279) /sn:0 /w:[ 0 ]

endmodule

module CSA_4bit(S, Co, B, Ci, A);
//: interface  /sz:(156, 142) /bd:[ Ti0>B[3:0](169/254) Ti1>A[3:0](72/254) Ri0>Ci(106/208) Lo0<Co(105/208) Bo0<S[3:0](123/254) ]
input [3:0] B;    //: /sn:0 {0}(778,382)(778,321)(596,321)(596,98){1}
//: {2}(598,96)(773,96)(773,135){3}
//: {4}(594,96)(503,96){5}
input [3:0] A;    //: /sn:0 {0}(694,382)(694,342)(557,342)(557,67){1}
//: {2}(559,65)(688,65)(688,135){3}
//: {4}(555,65)(504,65){5}
supply1 w0;    //: /sn:0 /dp:1 {0}(831,438)(894,438)(894,416){1}
supply0 w1;    //: /sn:0 {0}(884,204)(884,187)(827,187){1}
output Co;    //: /sn:0 /dp:1 {0}(435,302)(393,302){1}
input Ci;    //: /sn:0 {0}(377,597)(404,597){1}
//: {2}(406,595)(406,573)(330,573)(330,245)(448,245)(448,279){3}
//: {4}(406,599)(406,650)(697,650){5}
output [3:0] S;    //: /sn:0 {0}(720,709)(720,663){1}
wire [3:0] w6;    //: /sn:0 /dp:1 {0}(710,634)(710,596)(938,596)(938,307)(725,307)(725,276){1}
wire w7;    //: /sn:0 {0}(637,497)(476,497)(476,312)(464,312){1}
wire [3:0] w14;    //: /sn:0 {0}(730,634)(730,534){1}
wire w5;    //: /sn:0 {0}(630,242)(474,242)(474,292)(464,292){1}
//: enddecls

  //: output g4 (S) @(720,706) /sn:0 /R:3 /w:[ 0 ]
  //: joint g8 (A) @(557, 65) /w:[ 2 -1 4 1 ]
  //: output g3 (Co) @(396,302) /sn:0 /R:2 /w:[ 1 ]
  //: supply1 g2 (w0) @(905,416) /sn:0 /w:[ 1 ]
  //: input g1 (B) @(501,96) /sn:0 /w:[ 5 ]
  mux g10 (.I0(w5), .I1(w7), .S(Ci), .Z(Co));   //: @(448,302) /sn:0 /R:3 /w:[ 1 1 3 0 ] /ss:0 /do:0
  CPA g6 (.A(A), .B(B), .Ci(w1), .Co(w5), .S(w6));   //: @(631, 136) /sz:(195, 139) /sn:0 /p:[ Ti0>3 Ti1>3 Ri0>1 Lo0<0 Bo0<1 ]
  CPA g7 (.A(A), .B(B), .Ci(w0), .Co(w7), .S(w14));   //: @(638, 383) /sz:(192, 150) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>0 Lo0<0 Bo0<1 ]
  //: joint g9 (B) @(596, 96) /w:[ 2 -1 4 1 ]
  mux g12 (.I0(w6), .I1(w14), .S(Ci), .Z(S));   //: @(720,650) /sn:0 /w:[ 0 0 5 1 ] /ss:0 /do:0
  //: input g11 (Ci) @(375,597) /sn:0 /w:[ 0 ]
  //: supply0 g5 (w1) @(884,210) /sn:0 /w:[ 0 ]
  //: input g0 (A) @(502,65) /sn:0 /w:[ 5 ]
  //: joint g13 (Ci) @(406, 597) /w:[ -1 2 1 4 ]

endmodule

module CPA(B, Ci, Co, S, A);
//: interface  /sz:(190, 97) /bd:[ Ti0>A[3:0](56/190) Ti1>B[3:0](139/190) Ri0>Ci(36/97) Lo0<Co(74/97) Bo0<S[3:0](92/190) ]
input [3:0] B;    //: /sn:0 {0}(147,91)(246,91){1}
//: {2}(247,91)(544,91){3}
//: {4}(545,91)(825,91){5}
//: {6}(826,91)(1100,91){7}
//: {8}(1101,91)(1125,91){9}
input [3:0] A;    //: /sn:0 /dp:9 {0}(1086,156)(1051,156){1}
//: {2}(1050,156)(776,156){3}
//: {4}(775,156)(494,156){5}
//: {6}(493,156)(196,156){7}
//: {8}(195,156)(150,156){9}
output Co;    //: /sn:0 /dp:1 {0}(1128,328)(1228,328){1}
input Ci;    //: /sn:0 {0}(124,340)(166,340){1}
output [3:0] S;    //: /sn:0 /dp:1 {0}(1170,494)(1284,494){1}
wire w16;    //: /sn:0 {0}(572,334)(746,334){1}
wire w13;    //: /sn:0 {0}(513,382)(513,499)(1164,499){1}
wire w6;    //: /sn:0 {0}(1051,160)(1051,264)(1050,264)(1050,274){1}
wire w7;    //: /sn:0 {0}(1101,95)(1101,274){1}
wire w4;    //: /sn:0 {0}(196,160)(196,283){1}
wire w22;    //: /sn:0 {0}(854,331)(1020,331){1}
wire w3;    //: /sn:0 {0}(826,95)(826,267)(827,267)(827,277){1}
wire w0;    //: /sn:0 {0}(494,160)(494,280){1}
wire w20;    //: /sn:0 {0}(1164,489)(795,489)(795,379){1}
wire w1;    //: /sn:0 {0}(776,160)(776,277){1}
wire w27;    //: /sn:0 {0}(1164,479)(1069,479)(1069,376){1}
wire w14;    //: /sn:0 {0}(274,337)(464,337){1}
wire w2;    //: /sn:0 {0}(545,95)(545,280){1}
wire w15;    //: /sn:0 {0}(215,385)(215,509)(1164,509){1}
wire w5;    //: /sn:0 {0}(247,95)(247,283){1}
//: enddecls

  //: input g4 (B) @(145,91) /sn:0 /w:[ 0 ]
  tran g16(.Z(w4), .I(A[0]));   //: @(196,154) /sn:0 /R:1 /w:[ 0 8 7 ] /ss:1
  //: input g3 (Ci) @(122,340) /sn:0 /w:[ 0 ]
  tran g17(.Z(w2), .I(B[1]));   //: @(545,89) /sn:0 /R:1 /w:[ 0 3 4 ] /ss:1
  FA g2 (.B(w3), .A(w1), .Ci(w16), .S(w20), .Co(w22));   //: @(747, 278) /sz:(106, 100) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>1 Bo0<1 Ro0<0 ]
  //: output g23 (Co) @(1225,328) /sn:0 /w:[ 1 ]
  FA g1 (.B(w2), .A(w0), .Ci(w14), .S(w13), .Co(w16));   //: @(465, 281) /sz:(106, 100) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>1 Bo0<0 Ro0<0 ]
  //: output g24 (S) @(1281,494) /sn:0 /w:[ 1 ]
  tran g18(.Z(w0), .I(A[1]));   //: @(494,154) /sn:0 /R:1 /w:[ 0 6 5 ] /ss:1
  concat g25 (.I0(w15), .I1(w13), .I2(w20), .I3(w27), .Z(S));   //: @(1169,494) /sn:0 /w:[ 1 1 0 0 0 ] /dr:0
  FA g6 (.B(w7), .A(w6), .Ci(w22), .S(w27), .Co(Co));   //: @(1021, 275) /sz:(106, 100) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>1 Bo0<1 Ro0<0 ]
  tran g22(.Z(w6), .I(A[3]));   //: @(1051,154) /sn:0 /R:1 /w:[ 0 2 1 ] /ss:1
  //: input g5 (A) @(148,156) /sn:0 /w:[ 9 ]
  tran g21(.Z(w7), .I(B[3]));   //: @(1101,89) /sn:0 /R:1 /w:[ 0 7 8 ] /ss:1
  tran g19(.Z(w1), .I(A[2]));   //: @(776,154) /sn:0 /R:1 /w:[ 0 4 3 ] /ss:1
  tran g20(.Z(w3), .I(B[2]));   //: @(826,89) /sn:0 /R:1 /w:[ 0 5 6 ] /ss:1
  FA g0 (.B(w5), .A(w4), .Ci(Ci), .S(w15), .Co(w14));   //: @(167, 284) /sz:(106, 100) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>1 Bo0<0 Ro0<0 ]
  tran g15(.Z(w5), .I(B[0]));   //: @(247,89) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:1

endmodule

module FA(B, A, S, Co, Ci);
//: interface  /sz:(106, 100) /bd:[ Ti0>A(29/106) Ti1>B(80/106) Li0>Ci(56/100) Bo0<S(48/106) Ro0<Co(53/100) ]
input B;    //: /sn:0 {0}(337,288)(441,288){1}
input A;    //: /sn:0 {0}(336,221)(441,221){1}
output Co;    //: /sn:0 /dp:1 {0}(1026,295)(1073,295){1}
input Ci;    //: /sn:0 {0}(706,291)(771,291){1}
output S;    //: /sn:0 /dp:1 {0}(921,227)(1078,227){1}
wire w3;    //: /sn:0 {0}(591,224)(771,224){1}
wire w8;    //: /sn:0 /dp:1 {0}(1005,292)(921,292){1}
wire w2;    //: /sn:0 {0}(591,289)(640,289)(640,332)(977,332)(977,297)(1005,297){1}
//: enddecls

  //: input g4 (B) @(335,288) /sn:0 /w:[ 0 ]
  //: input g3 (A) @(334,221) /sn:0 /w:[ 0 ]
  or g2 (.I0(w8), .I1(w2), .Z(Co));   //: @(1016,295) /sn:0 /delay:" 5" /w:[ 0 1 0 ]
  HA g1 (.A(w3), .B(Ci), .S(S), .C(w8));   //: @(772, 189) /sz:(148, 128) /sn:0 /p:[ Li0>1 Li1>1 Ro0<0 Ro1<1 ]
  //: output g6 (S) @(1075,227) /sn:0 /w:[ 1 ]
  //: output g7 (Co) @(1070,295) /sn:0 /w:[ 1 ]
  //: input g5 (Ci) @(704,291) /sn:0 /w:[ 0 ]
  HA g0 (.A(A), .B(B), .S(w3), .C(w2));   //: @(442, 186) /sz:(148, 128) /sn:0 /p:[ Li0>1 Li1>1 Ro0<0 Ro1<0 ]

endmodule

module main;    //: root_module
wire [15:0] A0;    //: /sn:0 {0}(466,72)(466,121){1}
wire Co0;    //: /sn:0 {0}(368,185)(407,185){1}
wire w0;    //: /sn:0 {0}(4624,147)(4614,147){1}
wire w1;    //: /sn:0 {0}(23275,-10811)(23275,-10801){1}
wire w2;    //: /sn:0 {0}(678,177)(657,177)(657,182)(635,182){1}
wire [15:0] S;    //: /sn:0 {0}(510,314)(510,249){1}
wire [15:0] B0;    //: /sn:0 {0}(544,72)(544,121){1}
//: enddecls

  //: switch g4 (w0) @(4642,147) /sn:0 /R:2 /w:[ 0 ] /st:0
  led g3 (.I(S));   //: @(510,321) /sn:0 /R:2 /w:[ 0 ] /type:3
  //: dip g2 (B0) @(544,62) /sn:0 /w:[ 0 ] /st:15
  //: dip g1 (A0) @(466,62) /sn:0 /w:[ 0 ] /st:4
  //: switch g6 (w2) @(696,177) /sn:0 /R:2 /w:[ 0 ] /st:0
  led g7 (.I(Co0));   //: @(361,185) /sn:0 /R:1 /w:[ 0 ] /type:3
  //: switch g5 (w1) @(23275,-10824) /sn:0 /R:3 /w:[ 0 ] /st:0
  CSA_16b g0 (.B(B0), .A(A0), .Cin(w2), .Co(Co0), .S(S));   //: @(408, 122) /sz:(226, 126) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<1 Bo0<1 ]

endmodule
