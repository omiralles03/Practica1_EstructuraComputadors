//: version "1.8.7"

module main;    //: root_module
wire w6;    //: /sn:0 {0}(296,73)(296,132){1}
wire w4;    //: /sn:0 {0}(327,162)(405,162){1}
wire w0;    //: /sn:0 {0}(175,175)(225,175){1}
wire w3;    //: /sn:0 {0}(327,201)(405,201){1}
wire w5;    //: /sn:0 {0}(253,73)(253,132){1}
//: enddecls

  led g4 (.I(w4));   //: @(412,162) /sn:0 /R:3 /w:[ 1 ] /type:2
  //: switch g3 (w0) @(158,175) /sn:0 /w:[ 0 ] /st:1
  //: switch g2 (w6) @(296,60) /sn:0 /R:3 /w:[ 0 ] /st:1
  //: switch g1 (w5) @(253,60) /sn:0 /R:3 /w:[ 0 ] /st:1
  led g5 (.I(w3));   //: @(412,201) /sn:0 /R:3 /w:[ 1 ] /type:2
  FA g0 (.A(w5), .B(w6), .Cin(w0), .Cout(w4), .S(w3));   //: @(226, 133) /sz:(100, 89) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>1 Ro0<0 Ro1<0 ]

endmodule

module FA(Cout, S, Cin, B, A);
//: interface  /sz:(100, 89) /bd:[ Ti0>A(27/100) Ti1>B(70/100) Li0>Cin(42/89) Ro0<Cout(29/89) Ro1<S(68/89) ]
input B;    //: /sn:0 {0}(398,307)(450,307){1}
//: {2}(454,307)(504,307){3}
//: {4}(452,309)(452,352)(556,352){5}
input A;    //: /sn:0 {0}(556,357)(438,357)(438,284){1}
//: {2}(440,282)(490,282)(490,302)(504,302){3}
//: {4}(436,282)(398,282){5}
input Cin;    //: /sn:0 {0}(398,321)(549,321){1}
//: {2}(551,319)(551,310)(560,310){3}
//: {4}(551,323)(551,332)(556,332){5}
output Cout;    //: /sn:0 /dp:1 {0}(626,344)(659,344){1}
output S;    //: /sn:0 /dp:1 {0}(581,308)(659,308){1}
wire w14;    //: /sn:0 {0}(577,355)(596,355)(596,346)(605,346){1}
wire w2;    //: /sn:0 {0}(525,305)(537,305){1}
//: {2}(541,305)(560,305){3}
//: {4}(539,307)(539,337)(556,337){5}
wire w11;    //: /sn:0 {0}(577,335)(596,335)(596,341)(605,341){1}
//: enddecls

  //: output g4 (Cout) @(656,344) /sn:0 /w:[ 1 ]
  and g8 (.I0(Cin), .I1(w2), .Z(w11));   //: @(567,335) /sn:0 /delay:" 3" /w:[ 5 5 0 ]
  //: output g3 (S) @(656,308) /sn:0 /w:[ 1 ]
  //: input g2 (Cin) @(396,321) /sn:0 /w:[ 0 ]
  //: input g1 (B) @(396,307) /sn:0 /w:[ 0 ]
  //: joint g10 (Cin) @(551, 321) /w:[ -1 2 1 4 ]
  xor g6 (.I0(w2), .I1(Cin), .Z(S));   //: @(571,308) /sn:0 /delay:" 4" /w:[ 3 3 0 ]
  or g7 (.I0(w11), .I1(w14), .Z(Cout));   //: @(616,344) /sn:0 /delay:" 3" /w:[ 1 1 0 ]
  and g9 (.I0(B), .I1(A), .Z(w14));   //: @(567,355) /sn:0 /delay:" 3" /w:[ 5 0 0 ]
  //: joint g12 (B) @(452, 307) /w:[ 2 -1 1 4 ]
  //: joint g11 (A) @(438, 282) /w:[ 2 -1 4 1 ]
  xor g5 (.I0(A), .I1(B), .Z(w2));   //: @(515,305) /sn:0 /delay:" 4" /w:[ 3 3 0 ]
  //: input g0 (A) @(396,282) /sn:0 /w:[ 5 ]
  //: joint g13 (w2) @(539, 305) /w:[ 2 -1 1 4 ]

endmodule
