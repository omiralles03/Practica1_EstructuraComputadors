//: version "1.8.7"

module HA(C, S, B, A);
//: interface  /sz:(97, 93) /bd:[ Li0>A(25/93) Li1>B(65/93) Ro0<S(25/93) Ro1<C(66/93) ]
input B;    //: /sn:0 {0}(229,171)(256,171){1}
//: {2}(260,171)(287,171){3}
//: {4}(258,173)(258,197)(287,197){5}
input A;    //: /sn:0 {0}(228,146)(243,146)(243,166)(272,166){1}
//: {2}(276,166)(287,166){3}
//: {4}(274,168)(274,192)(287,192){5}
output C;    //: /sn:0 /dp:1 {0}(308,195)(341,195){1}
output S;    //: /sn:0 /dp:1 {0}(308,169)(340,169){1}
//: enddecls

  xor g4 (.I0(A), .I1(B), .Z(S));   //: @(298,169) /sn:0 /delay:" 4" /w:[ 3 3 0 ]
  //: output g3 (C) @(338,195) /sn:0 /w:[ 1 ]
  //: output g2 (S) @(337,169) /sn:0 /w:[ 1 ]
  //: input g1 (B) @(227,171) /sn:0 /w:[ 0 ]
  //: joint g6 (A) @(274, 166) /w:[ 2 -1 1 4 ]
  //: joint g7 (B) @(258, 171) /w:[ 2 -1 1 4 ]
  and g5 (.I0(A), .I1(B), .Z(C));   //: @(298,195) /sn:0 /delay:" 3" /w:[ 5 5 0 ]
  //: input g0 (A) @(226,146) /sn:0 /w:[ 0 ]

endmodule

module main;    //: root_module
wire w6;    //: /sn:0 {0}(296,73)(296,132){1}
wire w4;    //: /sn:0 {0}(327,162)(405,162){1}
wire w0;    //: /sn:0 {0}(175,175)(225,175){1}
wire w3;    //: /sn:0 {0}(327,201)(405,201){1}
wire w5;    //: /sn:0 {0}(253,73)(253,132){1}
//: enddecls

  led g4 (.I(w4));   //: @(412,162) /sn:0 /R:3 /w:[ 1 ] /type:2
  //: switch g3 (w0) @(158,175) /sn:0 /w:[ 0 ] /st:1
  //: switch g2 (w6) @(296,60) /sn:0 /R:3 /w:[ 0 ] /st:1
  //: switch g1 (w5) @(253,60) /sn:0 /R:3 /w:[ 0 ] /st:1
  led g5 (.I(w3));   //: @(412,201) /sn:0 /R:3 /w:[ 1 ] /type:2
  FA g0 (.A(w5), .B(w6), .Cin(w0), .Cout(w4), .S(w3));   //: @(226, 133) /sz:(100, 89) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>1 Ro0<0 Ro1<0 ]

endmodule

module FA(Cout, S, Cin, B, A);
//: interface  /sz:(100, 89) /bd:[ Ti0>A(27/100) Ti1>B(70/100) Li0>Cin(42/89) Ro0<Cout(29/89) Ro1<S(68/89) ]
input B;    //: /sn:0 {0}(413,322)(511,322){1}
input A;    //: /sn:0 {0}(409,282)(511,282){1}
input Cin;    //: /sn:0 {0}(407,238)(670,238){1}
output Cout;    //: /sn:0 {0}(871,287)(826,287){1}
output S;    //: /sn:0 /dp:1 {0}(769,243)(873,243){1}
wire w0;    //: /sn:0 /dp:1 {0}(805,284)(769,284){1}
wire w3;    //: /sn:0 {0}(610,323)(796,323)(796,289)(805,289){1}
wire w2;    //: /sn:0 {0}(610,282)(670,282){1}
//: enddecls

  //: output g4 (Cout) @(868,287) /sn:0 /w:[ 0 ]
  //: output g3 (S) @(870,243) /sn:0 /w:[ 1 ]
  //: input g2 (Cin) @(405,238) /sn:0 /w:[ 0 ]
  //: input g1 (B) @(411,322) /sn:0 /w:[ 0 ]
  HA g6 (.B(Cin), .A(w2), .C(w0), .S(S));   //: @(671, 218) /sz:(97, 93) /sn:0 /p:[ Li0>1 Li1>1 Ro0<1 Ro1<0 ]
  or g7 (.I0(w0), .I1(w3), .Z(Cout));   //: @(816,287) /sn:0 /delay:" 3" /w:[ 0 1 1 ]
  HA g5 (.B(B), .A(A), .C(w3), .S(w2));   //: @(512, 257) /sz:(97, 93) /sn:0 /p:[ Li0>1 Li1>1 Ro0<0 Ro1<0 ]
  //: input g0 (A) @(407,282) /sn:0 /w:[ 0 ]

endmodule
