//: version "1.8.7"

module CLL(Ci, C0, Pg, C4, G, P, Gg);
//: interface  /sz:(550, 62) /bd:[ Ti0>P[3:0](250/550) Ti1>G[3:0](125/550) Li0>C0(32/62) To0<Ci[2:0](384/550) Bo0<Pg(421/550) Bo1<Gg(477/550) Ro0<C4(30/62) ]
input C0;    //: /sn:0 {0}(326,481)(412,481){1}
input [3:0] G;    //: /sn:0 {0}(388,209)(491,209){1}
//: {2}(492,209)(649,209){3}
//: {4}(650,209)(816,209){5}
//: {6}(817,209)(986,209){7}
//: {8}(987,209)(1060,209){9}
output Pg;    //: /sn:0 /dp:1 {0}(964,86)(1009,86){1}
output C4;    //: /sn:0 {0}(1018,484)(1101,484){1}
input [3:0] P;    //: /sn:0 {0}(389,159)(448,159){1}
//: {2}(449,159)(606,159){3}
//: {4}(607,159)(773,159){5}
//: {6}(774,159)(943,159){7}
//: {8}(944,159)(1050,159){9}
output Gg;    //: /sn:0 /dp:1 {0}(1313,242)(1345,242){1}
input [2:0] Ci;    //: /sn:0 /dp:1 {0}(958,587)(989,587){1}
wire w6;    //: /sn:0 {0}(1114,253)(1131,253)(1131,240)(1292,240){1}
wire w13;    //: /sn:0 {0}(943,94)(886,94)(886,185)(942,185){1}
//: {2}(944,183)(944,163){3}
//: {4}(944,187)(944,248){5}
//: {6}(946,250)(1093,250){7}
//: {8}(944,252)(944,308){9}
//: {10}(946,310)(1093,310){11}
//: {12}(944,312)(944,352){13}
//: {14}(946,354)(1096,354){15}
//: {16}(944,356)(944,429){17}
wire w16;    //: /sn:0 /dp:1 {0}(848,484)(876,484){1}
//: {2}(880,484)(907,484){3}
//: {4}(878,486)(878,577)(952,577){5}
wire w4;    //: /sn:0 {0}(1096,364)(609,364){1}
//: {2}(607,362)(607,193){3}
//: {4}(609,191)(659,191)(659,84)(943,84){5}
//: {6}(607,189)(607,163){7}
//: {8}(607,366)(607,429){9}
wire w3;    //: /sn:0 {0}(1093,320)(652,320){1}
//: {2}(650,318)(650,213){3}
//: {4}(650,322)(650,429){5}
wire w0;    //: /sn:0 {0}(449,163)(449,184){1}
//: {2}(451,186)(535,186)(535,79)(943,79){3}
//: {4}(449,188)(449,426){5}
wire w12;    //: /sn:0 {0}(987,213)(987,233){1}
//: {2}(989,235)(1292,235){3}
//: {4}(987,237)(987,429){5}
wire w10;    //: /sn:0 {0}(570,481)(549,481){1}
//: {2}(545,481)(523,481){3}
//: {4}(547,483)(547,597)(952,597){5}
wire w1;    //: /sn:0 {0}(1292,245)(1174,245)(1174,315)(1114,315){1}
wire w8;    //: /sn:0 {0}(817,213)(817,253){1}
//: {2}(819,255)(1093,255){3}
//: {4}(817,257)(817,429){5}
wire w17;    //: /sn:0 /dp:1 {0}(681,484)(705,484){1}
//: {2}(709,484)(737,484){3}
//: {4}(707,486)(707,587)(952,587){5}
wire w2;    //: /sn:0 {0}(1292,250)(1210,250)(1210,361)(1117,361){1}
wire w5;    //: /sn:0 {0}(1096,369)(494,369){1}
//: {2}(492,367)(492,213){3}
//: {4}(492,371)(492,426){5}
wire w9;    //: /sn:0 {0}(943,89)(827,89)(827,188)(776,188){1}
//: {2}(774,186)(774,163){3}
//: {4}(774,190)(774,313){5}
//: {6}(776,315)(1093,315){7}
//: {8}(774,317)(774,357){9}
//: {10}(776,359)(1096,359){11}
//: {12}(774,361)(774,429){13}
//: enddecls

  //: input g4 (Ci) @(991,587) /sn:0 /R:2 /w:[ 1 ]
  Ci g8 (.G(w8), .P(w9), .Ci(w17), .CO(w16));   //: @(738, 430) /sz:(109, 98) /sn:0 /p:[ Ti0>5 Ti1>13 Li0>3 Ro0<0 ]
  //: input g3 (C0) @(324,481) /sn:0 /w:[ 0 ]
  concat g16 (.I0(w10), .I1(w17), .I2(w16), .Z(Ci));   //: @(957,587) /sn:0 /w:[ 5 5 5 0 ] /dr:0
  //: output g26 (Pg) @(1006,86) /sn:0 /w:[ 1 ]
  //: output g17 (C4) @(1098,484) /sn:0 /w:[ 1 ]
  //: input g2 (G) @(386,209) /sn:0 /w:[ 0 ]
  or g30 (.I0(w12), .I1(w6), .I2(w1), .I3(w2), .Z(Gg));   //: @(1303,242) /sn:0 /delay:" 5" /w:[ 3 1 0 0 0 ]
  //: joint g23 (w4) @(607, 191) /w:[ 4 6 -1 3 ]
  //: joint g39 (w4) @(607, 364) /w:[ 1 2 -1 8 ]
  //: joint g24 (w9) @(774, 188) /w:[ 1 2 -1 4 ]
  //: input g1 (P) @(387,159) /sn:0 /w:[ 0 ]
  and g29 (.I0(w13), .I1(w9), .I2(w4), .I3(w5), .Z(w2));   //: @(1107,361) /sn:0 /delay:" 5" /w:[ 15 11 0 0 1 ]
  //: joint g18 (w10) @(547, 481) /w:[ 1 -1 2 4 ]
  //: joint g25 (w13) @(944, 185) /w:[ -1 2 1 4 ]
  tran g10(.Z(w4), .I(P[1]));   //: @(607,157) /sn:0 /R:1 /w:[ 7 3 4 ] /ss:1
  tran g6(.Z(w5), .I(G[0]));   //: @(492,207) /sn:0 /R:1 /w:[ 3 1 2 ] /ss:1
  //: joint g35 (w9) @(774, 315) /w:[ 6 5 -1 8 ]
  Ci g7 (.G(w3), .P(w4), .Ci(w10), .CO(w17));   //: @(571, 430) /sz:(109, 98) /sn:0 /p:[ Ti0>5 Ti1>9 Li0>0 Ro0<0 ]
  Ci g9 (.G(w12), .P(w13), .Ci(w16), .CO(C4));   //: @(908, 430) /sz:(109, 98) /sn:0 /p:[ Ti0>5 Ti1>17 Li0>3 Ro0<0 ]
  //: joint g31 (w12) @(987, 235) /w:[ 2 1 -1 4 ]
  //: joint g22 (w0) @(449, 186) /w:[ 2 1 -1 4 ]
  //: output g41 (Gg) @(1342,242) /sn:0 /w:[ 1 ]
  //: joint g36 (w3) @(650, 320) /w:[ 1 2 -1 4 ]
  //: joint g33 (w8) @(817, 255) /w:[ 2 1 -1 4 ]
  //: joint g40 (w5) @(492, 369) /w:[ 1 2 -1 4 ]
  tran g12(.Z(w9), .I(P[2]));   //: @(774,157) /sn:0 /R:1 /w:[ 3 5 6 ] /ss:1
  //: joint g34 (w13) @(944, 310) /w:[ 10 9 -1 12 ]
  and g28 (.I0(w13), .I1(w9), .I2(w3), .Z(w1));   //: @(1104,315) /sn:0 /delay:" 5" /w:[ 11 7 0 1 ]
  tran g5(.Z(w0), .I(P[0]));   //: @(449,157) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:1
  tran g11(.Z(w3), .I(G[1]));   //: @(650,207) /sn:0 /R:1 /w:[ 3 3 4 ] /ss:1
  tran g14(.Z(w13), .I(P[3]));   //: @(944,157) /sn:0 /R:1 /w:[ 3 7 8 ] /ss:1
  and g21 (.I0(w0), .I1(w4), .I2(w9), .I3(w13), .Z(Pg));   //: @(954,86) /sn:0 /delay:" 5" /w:[ 3 5 0 0 0 ]
  //: joint g19 (w17) @(707, 484) /w:[ 2 -1 1 4 ]
  //: joint g32 (w13) @(944, 250) /w:[ 6 5 -1 8 ]
  //: joint g20 (w16) @(878, 484) /w:[ 2 -1 1 4 ]
  //: joint g38 (w9) @(774, 359) /w:[ 10 9 -1 12 ]
  Ci g0 (.G(w5), .P(w0), .Ci(C0), .CO(w10));   //: @(413, 427) /sz:(109, 99) /sn:0 /p:[ Ti0>5 Ti1>5 Li0>1 Ro0<3 ]
  tran g15(.Z(w12), .I(G[3]));   //: @(987,207) /sn:0 /R:1 /w:[ 0 7 8 ] /ss:1
  and g27 (.I0(w13), .I1(w8), .Z(w6));   //: @(1104,253) /sn:0 /delay:" 5" /w:[ 7 3 0 ]
  //: joint g37 (w13) @(944, 354) /w:[ 14 13 -1 16 ]
  tran g13(.Z(w8), .I(G[2]));   //: @(817,207) /sn:0 /R:1 /w:[ 0 5 6 ] /ss:1

endmodule

module PFA(B, S, A, Gi, Pi, Cin);
//: interface  /sz:(105, 86) /bd:[ Ti0>B(69/105) Ti1>A(35/105) Li0>Cin(41/86) Ro0<Pi(42/86) Ro1<Gi(64/86) Ro2<S(20/86) ]
input B;    //: /sn:0 {0}(312,108)(254,108){1}
//: {2}(250,108)(207,108){3}
//: {4}(252,110)(252,153){5}
//: {6}(254,155)(405,155){7}
//: {8}(252,157)(252,183)(404,183){9}
output Gi;    //: /sn:0 {0}(425,181)(453,181){1}
input A;    //: /sn:0 {0}(207,98)(281,98){1}
//: {2}(285,98)(302,98)(302,103)(312,103){3}
//: {4}(283,100)(283,148){5}
//: {6}(285,150)(405,150){7}
//: {8}(283,152)(283,178)(404,178){9}
input Cin;    //: /sn:0 {0}(199,136)(227,136)(227,127)(403,127){1}
output Pi;    //: /sn:0 /dp:1 {0}(426,153)(453,153){1}
output S;    //: /sn:0 /dp:1 {0}(424,125)(449,125){1}
wire w2;    //: /sn:0 {0}(333,106)(400,106)(400,122)(403,122){1}
//: enddecls

  //: joint g4 (A) @(283, 98) /w:[ 2 -1 1 4 ]
  //: input g8 (B) @(205,108) /sn:0 /w:[ 3 ]
  and g3 (.I0(A), .I1(B), .Z(Gi));   //: @(415,181) /sn:0 /delay:" 5" /w:[ 9 9 0 ]
  or g2 (.I0(A), .I1(B), .Z(Pi));   //: @(416,153) /sn:0 /delay:" 5" /w:[ 7 7 0 ]
  xor g1 (.I0(w2), .I1(Cin), .Z(S));   //: @(414,125) /sn:0 /delay:" 6" /w:[ 1 1 0 ]
  //: output g10 (S) @(446,125) /sn:0 /w:[ 1 ]
  //: joint g6 (B) @(252, 108) /w:[ 1 -1 2 4 ]
  //: joint g7 (B) @(252, 155) /w:[ 6 5 -1 8 ]
  //: input g9 (A) @(205,98) /sn:0 /w:[ 0 ]
  //: output g12 (Gi) @(450,181) /sn:0 /w:[ 1 ]
  //: joint g5 (A) @(283, 150) /w:[ 6 5 -1 8 ]
  //: output g11 (Pi) @(450,153) /sn:0 /w:[ 1 ]
  xor g0 (.I0(A), .I1(B), .Z(w2));   //: @(323,106) /sn:0 /delay:" 6" /w:[ 3 0 0 ]
  //: input g13 (Cin) @(197,136) /sn:0 /w:[ 0 ]

endmodule

module Ci(CO, Ci, G, P);
//: interface  /sz:(109, 99) /bd:[ Ti0>P(36/109) Ti1>G(79/109) Li0>Ci(54/99) Ro0<CO(54/99) ]
output CO;    //: /sn:0 {0}(708,266)(669,266){1}
input G;    //: /sn:0 /dp:1 {0}(648,263)(624,263)(624,241)(578,241){1}
input P;    //: /sn:0 {0}(512,278)(545,278)(545,295)(578,295){1}
input Ci;    //: /sn:0 /dp:1 {0}(578,300)(545,300)(545,316)(513,316){1}
wire Co;    //: /sn:0 /dp:1 {0}(599,298)(623,298)(623,268)(648,268){1}
//: enddecls

  and g4 (.I0(P), .I1(Ci), .Z(Co));   //: @(589,298) /sn:0 /delay:" 5" /w:[ 1 0 0 ]
  //: output g3 (CO) @(705,266) /sn:0 /w:[ 0 ]
  //: input g2 (Ci) @(511,316) /sn:0 /w:[ 1 ]
  //: input g1 (G) @(576,241) /sn:0 /w:[ 1 ]
  or g5 (.I0(G), .I1(Co), .Z(CO));   //: @(659,266) /sn:0 /delay:" 5" /w:[ 0 1 1 ]
  //: input g0 (P) @(510,278) /sn:0 /w:[ 0 ]

endmodule

module main;    //: root_module
wire [15:0] w6;    //: /sn:0 /dp:1 {0}(639,168)(639,246){1}
wire [15:0] w7;    //: /sn:0 /dp:1 {0}(728,169)(728,246){1}
wire w0;    //: /sn:0 {0}(732,459)(732,496){1}
wire w3;    //: /sn:0 {0}(821,352)(868,352){1}
wire [15:0] w1;    //: /sn:0 {0}(632,498)(632,459){1}
wire w2;    //: /sn:0 {0}(789,459)(789,497){1}
wire w5;    //: /sn:0 {0}(501,346)(558,346){1}
//: enddecls

  led g4 (.I(w3));   //: @(875,352) /sn:0 /R:3 /w:[ 1 ] /type:3
  //: dip g3 (w7) @(728,159) /sn:0 /w:[ 0 ] /st:10
  //: dip g2 (w6) @(639,158) /sn:0 /w:[ 0 ] /st:65535
  //: switch g1 (w5) @(484,346) /sn:0 /w:[ 0 ] /st:1
  led g6 (.I(w0));   //: @(732,503) /sn:0 /R:2 /w:[ 1 ] /type:3
  led g7 (.I(w2));   //: @(789,504) /sn:0 /R:2 /w:[ 1 ] /type:3
  led g5 (.I(w1));   //: @(632,505) /sn:0 /R:2 /w:[ 0 ] /type:3
  CLA_16bit g0 (.B(w7), .A(w6), .Ci(w5), .Gg(w2), .Pg(w0), .S(w1), .Co(w3));   //: @(559, 247) /sz:(261, 211) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>1 Bo0<0 Bo1<0 Bo2<1 Ro0<0 ]

endmodule

module CLA_4b(C4, S, B, Pg, Gg, A, C0);
//: interface  /sz:(101, 87) /bd:[ Ti0>B[3:0](71/101) Ti1>A[3:0](25/101) Li0>C0(37/87) Bo0<S(47/101) Ro0<C4(39/87) ]
input [3:0] B;    //: /sn:0 {0}(317,123)(401,123){1}
//: {2}(402,123)(591,123){3}
//: {4}(592,123)(775,123){5}
//: {6}(776,123)(962,123){7}
//: {8}(963,123)(1022,123){9}
input C0;    //: /sn:0 {0}(269,244)(296,244){1}
//: {2}(300,244)(332,244){3}
//: {4}(298,246)(298,509)(389,509){5}
input [3:0] A;    //: /sn:0 {0}(317,83)(367,83){1}
//: {2}(368,83)(557,83){3}
//: {4}(558,83)(741,83){5}
//: {6}(742,83)(928,83){7}
//: {8}(929,83)(1027,83){9}
output Pg;    //: /sn:0 {0}(845,540)(845,583)(865,583){1}
output C4;    //: /sn:0 {0}(941,507)(996,507){1}
output Gg;    //: /sn:0 {0}(893,540)(893,584)(923,584){1}
output [3:0] S;    //: /sn:0 /dp:1 {0}(1281,160)(1212,160){1}
wire w6;    //: /sn:0 {0}(742,199)(742,87){1}
wire w13;    //: /sn:0 {0}(963,196)(963,127){1}
wire w16;    //: /sn:0 {0}(1000,261)(1009,261)(1009,383)(530,383)(530,445){1}
wire w7;    //: /sn:0 {0}(776,199)(776,127){1}
wire [3:0] w34;    //: /sn:0 {0}(640,451)(640,476){1}
wire w4;    //: /sn:0 {0}(439,267)(461,267)(461,389)(500,389)(500,445){1}
wire w25;    //: /sn:0 /dp:1 {0}(1206,155)(639,155)(639,222)(629,222){1}
wire w0;    //: /sn:0 {0}(368,202)(368,87){1}
wire w3;    //: /sn:0 {0}(439,223)(459,223)(459,145)(1206,145){1}
wire w22;    //: /sn:0 {0}(629,266)(637,266)(637,341)(510,341)(510,445){1}
wire [3:0] w29;    //: /sn:0 /dp:1 {0}(515,451)(515,476){1}
wire w12;    //: /sn:0 {0}(929,196)(929,87){1}
wire w18;    //: /sn:0 {0}(558,201)(558,87){1}
wire w19;    //: /sn:0 {0}(592,201)(592,127){1}
wire w10;    //: /sn:0 {0}(813,264)(821,264)(821,353)(520,353)(520,445){1}
wire w23;    //: /sn:0 {0}(629,244)(645,244)(645,445){1}
wire w1;    //: /sn:0 {0}(402,202)(402,127){1}
wire w17;    //: /sn:0 {0}(1000,239)(1051,239)(1051,393)(625,393)(625,445){1}
wire w27;    //: /sn:0 {0}(1206,165)(833,165)(833,220)(813,220){1}
wire w28;    //: /sn:0 {0}(1206,175)(1030,175)(1030,217)(1000,217){1}
wire w14;    //: /sn:0 {0}(893,238)(872,238)(872,368)(764,368)(764,436){1}
wire w11;    //: /sn:0 {0}(813,242)(850,242)(850,404)(635,404)(635,445){1}
wire w2;    //: /sn:0 /dp:1 {0}(784,436)(784,309)(503,309)(503,243)(522,243){1}
wire [2:0] w15;    //: /sn:0 /dp:1 {0}(774,442)(774,476){1}
wire w5;    //: /sn:0 {0}(439,245)(485,245)(485,362)(655,362)(655,445){1}
wire w9;    //: /sn:0 /dp:1 {0}(774,436)(774,331)(692,331)(692,240)(706,240){1}
//: enddecls

  PFA g4 (.B(w7), .A(w6), .Cin(w9), .Pi(w11), .Gi(w10), .S(w27));   //: @(707, 200) /sz:(105, 86) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>1 Ro0<0 Ro1<0 Ro2<1 ]
  tran g8(.Z(w1), .I(B[0]));   //: @(402,121) /sn:0 /R:1 /w:[ 1 1 2 ] /ss:1
  CLL g3 (.P(w34), .G(w29), .C0(C0), .Ci(w15), .Gg(Gg), .Pg(Pg), .C4(C4));   //: @(390, 477) /sz:(550, 62) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>5 To0<1 Bo0<0 Bo1<0 Ro0<0 ]
  //: output g16 (C4) @(993,507) /sn:0 /w:[ 1 ]
  //: output g17 (S) @(1278,160) /sn:0 /w:[ 0 ]
  //: input g2 (B) @(315,123) /sn:0 /w:[ 0 ]
  //: output g23 (Pg) @(862,583) /sn:0 /w:[ 1 ]
  //: output g24 (Gg) @(920,584) /sn:0 /w:[ 1 ]
  //: input g1 (A) @(315,83) /sn:0 /w:[ 0 ]
  //: joint g18 (C0) @(298, 244) /w:[ 2 -1 1 4 ]
  tran g10(.Z(w19), .I(B[1]));   //: @(592,121) /sn:0 /R:1 /w:[ 1 3 4 ] /ss:1
  PFA g6 (.B(w19), .A(w18), .Cin(w2), .Pi(w23), .Gi(w22), .S(w25));   //: @(523, 202) /sz:(105, 86) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>1 Ro0<0 Ro1<0 Ro2<1 ]
  tran g7(.Z(w0), .I(A[0]));   //: @(368,81) /sn:0 /R:1 /w:[ 1 1 2 ] /ss:1
  tran g9(.Z(w18), .I(A[1]));   //: @(558,81) /sn:0 /R:1 /w:[ 1 3 4 ] /ss:1
  concat g22 (.I0(w3), .I1(w25), .I2(w27), .I3(w28), .Z(S));   //: @(1211,160) /sn:0 /w:[ 1 0 0 0 1 ] /dr:1
  tran g12(.Z(w7), .I(B[2]));   //: @(776,121) /sn:0 /R:1 /w:[ 1 5 6 ] /ss:1
  PFA g5 (.B(w13), .A(w12), .Cin(w14), .Pi(w17), .Gi(w16), .S(w28));   //: @(894, 197) /sz:(105, 86) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>0 Ro0<0 Ro1<0 Ro2<1 ]
  tran g11(.Z(w6), .I(A[2]));   //: @(742,81) /sn:0 /R:1 /w:[ 1 5 6 ] /ss:1
  tran g14(.Z(w13), .I(B[3]));   //: @(963,121) /sn:0 /R:1 /w:[ 1 7 8 ] /ss:1
  concat g19 (.I0(w4), .I1(w22), .I2(w10), .I3(w16), .Z(w29));   //: @(515,450) /sn:0 /R:3 /w:[ 1 1 1 1 0 ] /dr:0
  concat g21 (.I0(w2), .I1(w9), .I2(w14), .Z(w15));   //: @(774,441) /sn:0 /R:3 /w:[ 0 0 1 0 ] /dr:1
  concat g20 (.I0(w5), .I1(w23), .I2(w11), .I3(w17), .Z(w34));   //: @(640,450) /sn:0 /R:3 /w:[ 1 1 1 1 0 ] /dr:1
  PFA g0 (.B(w1), .A(w0), .Cin(C0), .Pi(w5), .Gi(w4), .S(w3));   //: @(333, 203) /sz:(105, 86) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>3 Ro0<0 Ro1<0 Ro2<0 ]
  //: input g15 (C0) @(267,244) /sn:0 /w:[ 0 ]
  tran g13(.Z(w12), .I(A[3]));   //: @(929,81) /sn:0 /R:1 /w:[ 1 7 8 ] /ss:1

endmodule

module CLA_16bit(A, Co, Gg, B, Ci, S, Pg);
//: interface  /sz:(261, 211) /bd:[ Ti0>A[15:0](80/261) Ti1>B[15:0](169/261) Li0>Ci(99/211) Bo0<S[15:0](73/261) Bo1<Pg(173/261) Bo2<Gg(230/261) Ro0<Co(105/211) ]
input [15:0] B;    //: /sn:0 {0}(245,169)(438,169){1}
//: {2}(439,169)(618,169){3}
//: {4}(619,169)(795,169){5}
//: {6}(796,169)(973,169){7}
//: {8}(974,169)(1065,169){9}
input [15:0] A;    //: /sn:0 {0}(249,135)(392,135){1}
//: {2}(393,135)(572,135){3}
//: {4}(573,135)(749,135){5}
//: {6}(750,135)(927,135){7}
//: {8}(928,135)(1066,135){9}
output Pg;    //: /sn:0 {0}(816,586)(816,545){1}
output Co;    //: /sn:0 /dp:1 {0}(922,512)(999,512){1}
output Gg;    //: /sn:0 {0}(856,582)(856,545){1}
input Ci;    //: /sn:0 {0}(370,514)(324,514)(324,257){1}
//: {2}(326,255)(367,255){3}
//: {4}(322,255)(297,255){5}
output [15:0] S;    //: /sn:0 /dp:1 {0}(1198,641)(1253,641){1}
wire w13;    //: /sn:0 {0}(511,451)(511,412)(990,412)(990,309){1}
wire [3:0] w6;    //: /sn:0 {0}(619,218)(619,173){1}
wire [3:0] w16;    //: /sn:0 {0}(974,220)(974,173){1}
wire [3:0] w7;    //: /sn:0 {0}(657,456)(657,481){1}
wire w39;    //: /sn:0 {0}(662,450)(662,357)(793,357)(793,308){1}
wire [3:0] w25;    //: /sn:0 /dp:1 {0}(1192,656)(415,656)(415,306){1}
wire w4;    //: /sn:0 /dp:1 {0}(679,229)(679,258)(650,258){1}
wire w36;    //: /sn:0 /dp:1 {0}(968,309)(968,366)(672,366)(672,450){1}
wire w22;    //: /sn:0 {0}(864,456)(864,445)(878,445)(878,258)(902,258){1}
wire w3;    //: /sn:0 {0}(439,306)(439,354)(642,354)(642,450){1}
wire [3:0] w0;    //: /sn:0 {0}(393,217)(393,139){1}
wire w30;    //: /sn:0 /dp:1 {0}(844,456)(844,428)(533,428)(533,256)(547,256){1}
wire w12;    //: /sn:0 {0}(458,306)(458,417)(481,417)(481,451){1}
wire [3:0] w18;    //: /sn:0 /dp:1 {0}(941,309)(941,626)(1192,626){1}
wire [3:0] w10;    //: /sn:0 {0}(750,219)(750,139){1}
wire w24;    //: /sn:0 /dp:1 {0}(497,234)(497,257)(470,257){1}
wire w31;    //: /sn:0 /dp:1 {0}(854,456)(854,436)(699,436)(699,257)(724,257){1}
wire [3:0] w1;    //: /sn:0 {0}(439,217)(439,173){1}
wire [2:0] w32;    //: /sn:0 /dp:1 {0}(854,462)(854,481){1}
wire [3:0] w8;    //: /sn:0 /dp:1 {0}(575,307)(575,646)(1192,646){1}
wire w17;    //: /sn:0 {0}(610,307)(610,343)(652,343)(652,450){1}
wire [3:0] w27;    //: /sn:0 /dp:1 {0}(496,457)(496,481){1}
wire w35;    //: /sn:0 /dp:1 {0}(812,308)(812,401)(501,401)(501,451){1}
wire [3:0] w28;    //: /sn:0 /dp:1 {0}(1192,636)(772,636)(772,308){1}
wire w14;    //: /sn:0 /dp:1 {0}(1049,248)(1049,260)(1005,260){1}
wire [3:0] w11;    //: /sn:0 {0}(796,219)(796,173){1}
wire [3:0] w15;    //: /sn:0 {0}(928,220)(928,139){1}
wire [3:0] w5;    //: /sn:0 {0}(573,218)(573,139){1}
wire w26;    //: /sn:0 {0}(491,451)(491,392)(630,392)(630,307){1}
wire w9;    //: /sn:0 /dp:1 {0}(861,249)(861,259)(827,259){1}
//: enddecls

  //: input g4 (A) @(247,135) /sn:0 /w:[ 0 ]
  tran g8(.Z(w5), .I(A[7:4]));   //: @(573,133) /sn:0 /R:1 /w:[ 1 3 4 ] /ss:1
  led g16 (.I(w24));   //: @(497,227) /sn:0 /w:[ 0 ] /type:0
  CLA_4b g3 (.B(w16), .A(w15), .C0(w22), .Gg(w13), .Pg(w36), .S(w18), .C4(w14));   //: @(903, 221) /sz:(101, 87) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>1 Bo0<1 Bo1<0 Bo2<0 Ro0<1 ]
  concat g26 (.I0(w30), .I1(w31), .I2(w22), .Z(w32));   //: @(854,461) /sn:0 /R:3 /w:[ 0 0 0 0 ] /dr:0
  led g17 (.I(w4));   //: @(679,222) /sn:0 /w:[ 0 ] /type:0
  CLA_4b g2 (.B(w11), .A(w10), .C0(w31), .Gg(w35), .Pg(w39), .S(w28), .C4(w9));   //: @(725, 220) /sz:(101, 87) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>1 Bo0<0 Bo1<1 Bo2<1 Ro0<1 ]
  concat g23 (.I0(w12), .I1(w26), .I2(w35), .I3(w13), .Z(w27));   //: @(496,456) /sn:0 /R:3 /w:[ 1 0 1 0 0 ] /dr:0
  concat g24 (.I0(w3), .I1(w17), .I2(w39), .I3(w36), .Z(w7));   //: @(657,455) /sn:0 /R:3 /w:[ 1 1 0 1 0 ] /dr:0
  CLA_4b g1 (.B(w6), .A(w5), .C0(w30), .Gg(w26), .Pg(w17), .S(w8), .C4(w4));   //: @(548, 219) /sz:(101, 87) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>1 Bo0<1 Bo1<0 Bo2<0 Ro0<1 ]
  led g18 (.I(w9));   //: @(861,242) /sn:0 /w:[ 0 ] /type:0
  //: output g25 (Co) @(996,512) /sn:0 /w:[ 1 ]
  tran g10(.Z(w10), .I(A[11:8]));   //: @(750,133) /sn:0 /R:1 /w:[ 1 5 6 ] /ss:1
  tran g6(.Z(w0), .I(A[3:0]));   //: @(393,133) /sn:0 /R:1 /w:[ 1 1 2 ] /ss:1
  tran g7(.Z(w1), .I(B[3:0]));   //: @(439,167) /sn:0 /R:1 /w:[ 1 1 2 ] /ss:1
  tran g9(.Z(w6), .I(B[7:4]));   //: @(619,167) /sn:0 /R:1 /w:[ 1 3 4 ] /ss:1
  concat g22 (.I0(w25), .I1(w8), .I2(w28), .I3(w18), .Z(S));   //: @(1197,641) /sn:0 /w:[ 0 1 0 1 0 ] /dr:0
  tran g12(.Z(w15), .I(A[15:12]));   //: @(928,133) /sn:0 /R:1 /w:[ 1 7 8 ] /ss:1
  //: output g28 (Gg) @(856,579) /sn:0 /R:3 /w:[ 0 ]
  //: input g5 (B) @(243,169) /sn:0 /w:[ 0 ]
  tran g11(.Z(w11), .I(B[11:8]));   //: @(796,167) /sn:0 /R:1 /w:[ 1 5 6 ] /ss:1
  //: input g14 (Ci) @(295,255) /sn:0 /w:[ 5 ]
  //: output g21 (S) @(1250,641) /sn:0 /w:[ 1 ]
  led g19 (.I(w14));   //: @(1049,241) /sn:0 /w:[ 0 ] /type:0
  //: joint g20 (Ci) @(324, 255) /w:[ 2 -1 4 1 ]
  CLL g15 (.G(w27), .P(w7), .C0(Ci), .Ci(w32), .Gg(Gg), .Pg(Pg), .C4(Co));   //: @(371, 482) /sz:(550, 62) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>0 To0<1 Bo0<1 Bo1<1 Ro0<0 ]
  CLA_4b g0 (.B(w1), .A(w0), .C0(Ci), .Gg(w12), .Pg(w3), .S(w25), .C4(w24));   //: @(368, 218) /sz:(101, 87) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>3 Bo0<0 Bo1<0 Bo2<1 Ro0<1 ]
  //: output g27 (Pg) @(816,583) /sn:0 /R:3 /w:[ 0 ]
  tran g13(.Z(w16), .I(B[15:12]));   //: @(974,167) /sn:0 /R:1 /w:[ 1 7 8 ] /ss:1

endmodule
