//: version "1.8.7"

module HA(C, S, B, A);
//: interface  /sz:(71, 65) /bd:[ Ti0>B(21/71) Ti1>A(53/71) Lo0<C(49/90) Bo0<S(49/100) ]
input B;    //: /sn:0 {0}(229,171)(256,171){1}
//: {2}(260,171)(287,171){3}
//: {4}(258,173)(258,197)(287,197){5}
input A;    //: /sn:0 {0}(228,146)(243,146)(243,166)(272,166){1}
//: {2}(276,166)(287,166){3}
//: {4}(274,168)(274,192)(287,192){5}
output C;    //: /sn:0 /dp:1 {0}(308,195)(341,195){1}
output S;    //: /sn:0 /dp:1 {0}(308,169)(340,169){1}
//: enddecls

  xor g4 (.I0(A), .I1(B), .Z(S));   //: @(298,169) /sn:0 /delay:" 4" /w:[ 3 3 0 ]
  //: output g3 (C) @(338,195) /sn:0 /w:[ 1 ]
  //: output g2 (S) @(337,169) /sn:0 /w:[ 1 ]
  //: input g1 (B) @(227,171) /sn:0 /w:[ 0 ]
  //: joint g6 (A) @(274, 166) /w:[ 2 -1 1 4 ]
  //: joint g7 (B) @(258, 171) /w:[ 2 -1 1 4 ]
  and g5 (.I0(A), .I1(B), .Z(C));   //: @(298,195) /sn:0 /delay:" 3" /w:[ 5 5 0 ]
  //: input g0 (A) @(226,146) /sn:0 /w:[ 0 ]

endmodule

module RCA_4b(Z, Y, X);
//: interface  /sz:(108, 99) /bd:[ Ti0>X[3:0](30/108) Ti1>Y[3:0](76/108) Bo0<Z[7:0](55/108) ]
input [3:0] X;    //: /sn:0 {0}(1242,258)(1138,258){1}
//: {2}(1136,256)(1136,104)(1017,104){3}
//: {4}(1016,104)(930,104){5}
//: {6}(929,104)(897,104){7}
//: {8}(896,104)(813,104){9}
//: {10}(812,104)(788,104){11}
//: {12}(787,104)(692,104){13}
//: {14}(691,104)(667,104){15}
//: {16}(666,104)(573,104){17}
//: {18}(572,104)(567,104){19}
//: {20}(1136,260)(1136,304){21}
//: {22}(1134,306)(833,306){23}
//: {24}(832,306)(705,306){25}
//: {26}(704,306)(579,306){27}
//: {28}(578,306)(458,306){29}
//: {30}(457,306)(451,306){31}
//: {32}(1136,308)(1136,475)(725,475){33}
//: {34}(724,475)(592,475){35}
//: {36}(591,475)(471,475){37}
//: {38}(470,475)(354,475){39}
//: {40}(353,475)(347,475){41}
output [7:0] Z;    //: /sn:0 /dp:1 {0}(1238,634)(1271,634){1}
input [3:0] Y;    //: /sn:0 {0}(1221,318)(1240,318){1}
wire w16;    //: /sn:0 /dp:1 {0}(672,128)(672,87)(791,87){1}
//: {2}(795,87)(901,87){3}
//: {4}(905,87)(1020,87){5}
//: {6}(1024,87)(1173,87)(1173,303)(1215,303){7}
//: {8}(1022,89)(1022,127){9}
//: {10}(903,89)(903,126){11}
//: {12}(793,89)(793,126){13}
wire w13;    //: /sn:0 {0}(901,147)(901,218){1}
wire w6;    //: /sn:0 {0}(841,254)(879,254){1}
wire w65;    //: /sn:0 {0}(382,577)(425,577){1}
wire w7;    //: /sn:0 {0}(804,286)(804,379){1}
wire w34;    //: /sn:0 {0}(354,479)(354,511){1}
wire w50;    //: /sn:0 {0}(607,416)(659,416){1}
wire w59;    //: /sn:0 {0}(836,363)(836,379){1}
wire w4;    //: /sn:0 {0}(579,310)(579,345){1}
wire w62;    //: /sn:0 {0}(463,347)(463,323)(582,323){1}
//: {2}(586,323)(708,323){3}
//: {4}(712,323)(836,323){5}
//: {6}(840,323)(1215,323){7}
//: {8}(838,325)(838,342){9}
//: {10}(710,325)(710,341){11}
//: {12}(584,325)(584,345){13}
wire w39;    //: /sn:0 {0}(695,202)(695,220){1}
wire w56;    //: /sn:0 {0}(357,532)(357,542){1}
wire w3;    //: /sn:0 {0}(833,310)(833,342){1}
wire w0;    //: /sn:0 {0}(1017,108)(1017,127){1}
wire w36;    //: /sn:0 {0}(791,147)(791,219){1}
wire w60;    //: /sn:0 /dp:1 {0}(462,608)(462,649)(1232,649){1}
wire w20;    //: /sn:0 {0}(1232,629)(709,629)(709,606){1}
wire w30;    //: /sn:0 {0}(592,479)(592,509){1}
wire w29;    //: /sn:0 {0}(733,415)(782,415){1}
wire w37;    //: /sn:0 {0}(667,108)(667,128){1}
wire w42;    //: /sn:0 {0}(670,149)(670,220){1}
wire w12;    //: /sn:0 {0}(582,366)(582,381){1}
wire w18;    //: /sn:0 {0}(720,255)(767,255){1}
wire w19;    //: /sn:0 {0}(1232,619)(817,619)(817,446){1}
wire w10;    //: /sn:0 {0}(458,310)(458,347){1}
wire w63;    //: /sn:0 /dp:1 {0}(1215,333)(1162,333)(1162,492)(732,492){1}
//: {2}(728,492)(599,492){3}
//: {4}(595,492)(478,492){5}
//: {6}(474,492)(359,492)(359,511){7}
//: {8}(476,494)(476,509){9}
//: {10}(597,494)(597,509){11}
//: {12}(730,494)(730,507){13}
wire w23;    //: /sn:0 {0}(1232,659)(345,659)(345,609){1}
wire w54;    //: /sn:0 {0}(436,382)(436,257)(522,257){1}
wire w24;    //: /sn:0 {0}(1232,669)(287,669)(287,578)(308,578){1}
wire w21;    //: /sn:0 {0}(1232,639)(583,639)(583,607){1}
wire w1;    //: /sn:0 {0}(578,182)(578,162)(695,162){1}
//: {2}(699,162)(816,162){3}
//: {4}(820,162)(933,162){5}
//: {6}(937,162)(1160,162)(1160,313)(1215,313){7}
//: {8}(935,164)(935,186){9}
//: {10}(818,164)(818,182){11}
//: {12}(697,164)(697,181){13}
wire w31;    //: /sn:0 {0}(557,288)(557,381){1}
wire w32;    //: /sn:0 {0}(461,368)(461,382){1}
wire w53;    //: /sn:0 {0}(728,528)(728,539){1}
wire w46;    //: /sn:0 {0}(620,575)(674,575){1}
wire w8;    //: /sn:0 /dp:1 {0}(898,126)(898,108)(897,108)(897,108){1}
wire w52;    //: /sn:0 {0}(570,448)(570,540){1}
wire w44;    //: /sn:0 {0}(595,530)(595,540){1}
wire w27;    //: /sn:0 {0}(708,362)(708,380){1}
wire w17;    //: /sn:0 /dp:1 {0}(1232,609)(914,609)(914,285){1}
wire w35;    //: /sn:0 {0}(813,108)(813,182){1}
wire w28;    //: /sn:0 {0}(683,380)(683,287){1}
wire w33;    //: /sn:0 {0}(816,203)(816,219){1}
wire w69;    //: /sn:0 {0}(474,530)(474,541){1}
wire w45;    //: /sn:0 {0}(576,203)(576,221){1}
wire w14;    //: /sn:0 /dp:1 {0}(1232,599)(1020,599)(1020,148){1}
wire w2;    //: /sn:0 /dp:1 {0}(595,256)(646,256){1}
wire w11;    //: /sn:0 {0}(933,207)(933,218){1}
wire w47;    //: /sn:0 {0}(696,447)(696,539){1}
wire w15;    //: /sn:0 {0}(725,479)(725,507){1}
wire w5;    //: /sn:0 {0}(705,310)(705,341){1}
wire w38;    //: /sn:0 {0}(692,108)(692,181){1}
wire w55;    //: /sn:0 {0}(486,417)(533,417){1}
wire w43;    //: /sn:0 {0}(471,479)(471,509){1}
wire w64;    //: /sn:0 /dp:1 {0}(332,542)(332,418)(412,418){1}
wire w9;    //: /sn:0 /dp:1 {0}(788,126)(788,108){1}
wire w26;    //: /sn:0 {0}(930,108)(930,186){1}
wire w51;    //: /sn:0 {0}(499,576)(546,576){1}
wire w40;    //: /sn:0 {0}(573,108)(573,182){1}
wire w57;    //: /sn:0 {0}(449,449)(449,541){1}
//: enddecls

  //: joint g44 (w62) @(584, 323) /w:[ 2 -1 1 12 ]
  concat g8 (.I0(w16), .I1(w1), .I2(w62), .I3(w63), .Z(Y));   //: @(1220,318) /sn:0 /w:[ 7 7 7 0 0 ] /dr:1
  //: output g4 (Z) @(1268,634) /sn:0 /w:[ 1 ]
  HA g47 (.A(w53), .B(w47), .C(w46), .S(w20));   //: @(675, 540) /sz:(71, 65) /sn:0 /p:[ Ti0>1 Ti1>1 Lo0<1 Bo0<1 ]
  //: joint g16 (w1) @(935, 162) /w:[ 6 -1 5 8 ]
  FA g3 (.B(w36), .A(w33), .Cin(w6), .Cout(w18), .S(w7));   //: @(768, 220) /sz:(72, 65) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<1 Bo0<0 ]
  //: joint g26 (w1) @(818, 162) /w:[ 4 -1 3 10 ]
  and g17 (.I0(w35), .I1(w1), .Z(w33));   //: @(816,193) /sn:0 /R:3 /delay:" 3" /w:[ 1 11 0 ]
  HA g2 (.A(w11), .B(w13), .C(w6), .S(w17));   //: @(880, 219) /sz:(71, 65) /sn:0 /p:[ Ti0>1 Ti1>1 Lo0<1 Bo0<1 ]
  //: joint g30 (w62) @(838, 323) /w:[ 6 -1 5 8 ]
  tran g23(.Z(w26), .I(X[0]));   //: @(930,102) /sn:0 /R:1 /w:[ 0 6 5 ] /ss:1
  //: joint g24 (w16) @(903, 87) /w:[ 4 -1 3 10 ]
  //: input g1 (Y) @(1242,318) /sn:0 /R:2 /w:[ 1 ]
  and g39 (.I0(w5), .I1(w62), .Z(w27));   //: @(708,352) /sn:0 /R:3 /delay:" 3" /w:[ 1 11 0 ]
  tran g60(.Z(w43), .I(X[2]));   //: @(471,473) /sn:0 /R:1 /w:[ 0 38 37 ] /ss:1
  tran g29(.Z(w9), .I(X[2]));   //: @(788,102) /sn:0 /R:1 /w:[ 1 12 11 ] /ss:1
  //: joint g51 (w63) @(730, 492) /w:[ 1 -1 2 12 ]
  and g18 (.I0(w9), .I1(w16), .Z(w36));   //: @(791,137) /sn:0 /R:3 /delay:" 3" /w:[ 0 13 0 ]
  tran g25(.Z(w8), .I(X[1]));   //: @(897,102) /sn:0 /R:1 /w:[ 1 8 7 ] /ss:1
  concat g10 (.I0(w14), .I1(w17), .I2(w19), .I3(w20), .I4(w21), .I5(w60), .I6(w23), .I7(w24), .Z(Z));   //: @(1237,634) /sn:0 /w:[ 0 0 0 0 0 1 0 0 0 ] /dr:1
  FA g49 (.B(w52), .A(w44), .Cin(w46), .Cout(w51), .S(w21));   //: @(547, 541) /sz:(72, 65) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<1 Bo0<1 ]
  and g50 (.I0(w15), .I1(w63), .Z(w53));   //: @(728,518) /sn:0 /R:3 /delay:" 3" /w:[ 1 13 0 ]
  and g6 (.I0(w8), .I1(w16), .Z(w13));   //: @(901,137) /sn:0 /R:3 /delay:" 3" /w:[ 0 11 0 ]
  and g58 (.I0(w43), .I1(w63), .Z(w69));   //: @(474,520) /sn:0 /R:3 /delay:" 3" /w:[ 1 9 0 ]
  FA g56 (.B(w57), .A(w69), .Cin(w51), .Cout(w65), .S(w60));   //: @(426, 542) /sz:(72, 65) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<1 Bo0<0 ]
  //: joint g9 (w16) @(1022, 87) /w:[ 6 -1 5 8 ]
  FA g35 (.B(w54), .A(w32), .Cin(w55), .Cout(w64), .S(w57));   //: @(413, 383) /sz:(72, 65) /sn:0 /p:[ Ti0>0 Ti1>1 Ri0>0 Lo0<1 Bo0<0 ]
  and g7 (.I0(w0), .I1(w16), .Z(w14));   //: @(1020,138) /sn:0 /R:3 /delay:" 3" /w:[ 1 9 1 ]
  //: joint g59 (w63) @(476, 492) /w:[ 5 -1 6 8 ]
  tran g31(.Z(w37), .I(X[3]));   //: @(667,102) /sn:0 /R:1 /w:[ 0 16 15 ] /ss:1
  HA g22 (.A(w59), .B(w7), .C(w29), .S(w19));   //: @(783, 380) /sz:(71, 65) /sn:0 /p:[ Ti0>1 Ti1>1 Lo0<1 Bo0<1 ]
  //: joint g54 (w63) @(597, 492) /w:[ 3 -1 4 10 ]
  tran g45(.Z(w4), .I(X[2]));   //: @(579,304) /sn:0 /R:1 /w:[ 0 28 27 ] /ss:1
  tran g41(.Z(w5), .I(X[1]));   //: @(705,304) /sn:0 /R:1 /w:[ 0 26 25 ] /ss:1
  and g36 (.I0(w3), .I1(w62), .Z(w59));   //: @(836,353) /sn:0 /R:3 /delay:" 3" /w:[ 1 9 0 ]
  FA g33 (.B(w28), .A(w27), .Cin(w29), .Cout(w50), .S(w47));   //: @(660, 381) /sz:(72, 65) /sn:0 /p:[ Ti0>0 Ti1>1 Ri0>0 Lo0<1 Bo0<0 ]
  tran g52(.Z(w15), .I(X[0]));   //: @(725,473) /sn:0 /R:1 /w:[ 0 34 33 ] /ss:1
  //: joint g42 (w62) @(710, 323) /w:[ 4 -1 3 10 ]
  tran g40(.Z(w40), .I(X[3]));   //: @(573,102) /sn:0 /R:1 /w:[ 0 18 17 ] /ss:1
  HA g12 (.A(w45), .B(w2), .C(w54), .S(w31));   //: @(523, 222) /sz:(71, 65) /sn:0 /p:[ Ti0>1 Ri0>0 Lo0<1 Bo0<0 ]
  FA g57 (.B(w64), .A(w56), .Cin(w65), .Cout(w24), .S(w23));   //: @(309, 543) /sz:(72, 65) /sn:0 /p:[ Ti0>0 Ti1>1 Ri0>0 Lo0<1 Bo0<1 ]
  and g46 (.I0(w10), .I1(w62), .Z(w32));   //: @(461,358) /sn:0 /R:3 /delay:" 3" /w:[ 1 0 0 ]
  //: joint g28 (w16) @(793, 87) /w:[ 2 -1 1 12 ]
  FA g34 (.B(w31), .A(w12), .Cin(w50), .Cout(w55), .S(w52));   //: @(534, 382) /sz:(72, 65) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<1 Bo0<0 ]
  //: joint g14 (X) @(1136, 306) /w:[ -1 21 22 32 ]
  FA g11 (.B(w42), .A(w39), .Cin(w18), .Cout(w2), .S(w28));   //: @(647, 221) /sz:(72, 65) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<1 Bo0<1 ]
  and g5 (.I0(w26), .I1(w1), .Z(w11));   //: @(933,197) /sn:0 /R:3 /delay:" 3" /w:[ 1 9 0 ]
  and g61 (.I0(w34), .I1(w63), .Z(w56));   //: @(357,522) /sn:0 /R:3 /delay:" 3" /w:[ 1 7 0 ]
  and g21 (.I0(w40), .I1(w1), .Z(w45));   //: @(576,193) /sn:0 /R:3 /delay:" 3" /w:[ 1 0 0 ]
  and g19 (.I0(w38), .I1(w1), .Z(w39));   //: @(695,192) /sn:0 /R:3 /delay:" 3" /w:[ 1 13 0 ]
  //: joint g32 (w1) @(697, 162) /w:[ 2 -1 1 12 ]
  and g20 (.I0(w37), .I1(w16), .Z(w42));   //: @(670,139) /sn:0 /R:3 /delay:" 3" /w:[ 1 0 0 ]
  and g43 (.I0(w4), .I1(w62), .Z(w12));   //: @(582,356) /sn:0 /R:3 /delay:" 3" /w:[ 1 13 0 ]
  tran g38(.Z(w3), .I(X[0]));   //: @(833,304) /sn:0 /R:1 /w:[ 0 24 23 ] /ss:1
  tran g15(.Z(w0), .I(X[0]));   //: @(1017,102) /sn:0 /R:1 /w:[ 0 4 3 ] /ss:1
  //: input g0 (X) @(1244,258) /sn:0 /R:2 /w:[ 0 ]
  tran g48(.Z(w10), .I(X[3]));   //: @(458,304) /sn:0 /R:1 /w:[ 0 30 29 ] /ss:1
  tran g27(.Z(w35), .I(X[1]));   //: @(813,102) /sn:0 /R:1 /w:[ 0 10 9 ] /ss:1
  tran g62(.Z(w34), .I(X[3]));   //: @(354,473) /sn:0 /R:1 /w:[ 0 40 39 ] /ss:1
  tran g37(.Z(w38), .I(X[2]));   //: @(692,102) /sn:0 /R:1 /w:[ 0 14 13 ] /ss:1
  tran g55(.Z(w30), .I(X[1]));   //: @(592,473) /sn:0 /R:1 /w:[ 0 36 35 ] /ss:1
  and g53 (.I0(w30), .I1(w63), .Z(w44));   //: @(595,520) /sn:0 /R:3 /delay:" 3" /w:[ 1 11 0 ]
  //: joint g13 (X) @(1136, 258) /w:[ 1 2 -1 20 ]

endmodule

module FA(Cout, S, Cin, B, A);
//: interface  /sz:(72, 65) /bd:[ Ti0>A(68/100) Ti1>B(33/100) Ri0>Cin(48/91) Lo0<Cout(50/91) Bo0<S(50/100) ]
input B;    //: /sn:0 {0}(413,322)(511,322){1}
input A;    //: /sn:0 {0}(409,282)(511,282){1}
input Cin;    //: /sn:0 {0}(407,238)(670,238){1}
output Cout;    //: /sn:0 {0}(871,287)(826,287){1}
output S;    //: /sn:0 /dp:1 {0}(769,243)(873,243){1}
wire w3;    //: /sn:0 {0}(610,323)(796,323)(796,289)(805,289){1}
wire w0;    //: /sn:0 /dp:1 {0}(805,284)(769,284){1}
wire w2;    //: /sn:0 {0}(610,282)(670,282){1}
//: enddecls

  //: output g4 (Cout) @(868,287) /sn:0 /w:[ 0 ]
  //: output g3 (S) @(870,243) /sn:0 /w:[ 1 ]
  //: input g2 (Cin) @(405,238) /sn:0 /w:[ 0 ]
  //: input g1 (B) @(411,322) /sn:0 /w:[ 0 ]
  HA g6 (.B(Cin), .A(w2), .C(w0), .S(S));   //: @(671, 218) /sz:(97, 93) /sn:0 /p:[ Li0>1 Li1>1 Ro0<1 Ro1<0 ]
  or g7 (.I0(w0), .I1(w3), .Z(Cout));   //: @(816,287) /sn:0 /delay:" 3" /w:[ 0 1 1 ]
  HA g5 (.B(B), .A(A), .C(w3), .S(w2));   //: @(512, 257) /sz:(97, 93) /sn:0 /p:[ Li0>1 Li1>1 Ro0<0 Ro1<0 ]
  //: input g0 (A) @(407,282) /sn:0 /w:[ 0 ]

endmodule

module main;    //: root_module
wire [3:0] w4;    //: /sn:0 {0}(276,138)(246,138)(246,164){1}
wire [7:0] w0;    //: /sn:0 {0}(225,287)(225,265){1}
wire [3:0] w3;    //: /sn:0 /dp:1 {0}(164,138)(200,138)(200,164){1}
//: enddecls

  led g3 (.I(w0));   //: @(225,294) /sn:0 /R:2 /w:[ 0 ] /type:2
  //: dip g2 (w4) @(314,138) /sn:0 /R:3 /w:[ 0 ] /st:2
  //: dip g1 (w3) @(126,138) /sn:0 /R:1 /w:[ 0 ] /st:10
  RCA_4b g0 (.Y(w4), .X(w3), .Z(w0));   //: @(170, 165) /sz:(108, 99) /sn:0 /p:[ Ti0>1 Ti1>1 Bo0<1 ]

endmodule
