//: version "1.8.7"

module FA(S, Co, Ci, B, A);
//: interface  /sz:(115, 101) /bd:[ Ti0>B(78/115) Ti1>A(34/115) Ri0>Ci(39/101) Lo0<Co(44/101) Bo0<S(47/115) ]
input B;    //: /sn:0 {0}(386,265)(414,265)(414,246)(447,246){1}
//: {2}(451,246)(474,246){3}
//: {4}(449,248)(449,320)(580,320){5}
input A;    //: /sn:0 {0}(388,240)(427,240){1}
//: {2}(431,240)(466,240)(466,241)(474,241){3}
//: {4}(429,242)(429,325)(580,325){5}
output Co;    //: /sn:0 /dp:1 {0}(607,256)(742,256)(742,214)(752,214){1}
input Ci;    //: /sn:0 {0}(388,283)(534,283)(534,278)(544,278){1}
//: {2}(546,276)(546,258)(586,258){3}
//: {4}(546,280)(546,294)(574,294){5}
output S;    //: /sn:0 {0}(757,318)(688,318)(688,315)(678,315){1}
wire w0;    //: /sn:0 /dp:1 {0}(586,253)(540,253)(540,244)(518,244){1}
//: {2}(514,244)(495,244){3}
//: {4}(516,246)(516,299)(574,299){5}
wire w8;    //: /sn:0 {0}(595,297)(647,297)(647,312)(657,312){1}
wire w11;    //: /sn:0 {0}(601,323)(647,323)(647,317)(657,317){1}
//: enddecls

  and g8 (.I0(B), .I1(A), .Z(w11));   //: @(591,323) /sn:0 /delay:" 5" /w:[ 5 5 0 ]
  //: output g4 (S) @(754,318) /sn:0 /w:[ 0 ]
  //: output g3 (Co) @(749,214) /sn:0 /w:[ 1 ]
  //: input g2 (Ci) @(386,283) /sn:0 /w:[ 0 ]
  //: input g1 (B) @(384,265) /sn:0 /w:[ 0 ]
  //: joint g10 (w0) @(516, 244) /w:[ 1 -1 2 4 ]
  xor g6 (.I0(A), .I1(B), .Z(w0));   //: @(485,244) /sn:0 /delay:" 6" /w:[ 3 3 3 ]
  or g9 (.I0(w8), .I1(w11), .Z(S));   //: @(668,315) /sn:0 /delay:" 5" /w:[ 1 1 1 ]
  and g7 (.I0(Ci), .I1(w0), .Z(w8));   //: @(585,297) /sn:0 /delay:" 5" /w:[ 5 5 0 ]
  //: joint g12 (A) @(429, 240) /w:[ 2 -1 1 4 ]
  //: joint g11 (Ci) @(546, 278) /w:[ -1 2 1 4 ]
  xor g5 (.I0(w0), .I1(Ci), .Z(Co));   //: @(597,256) /sn:0 /delay:" 6" /w:[ 0 3 0 ]
  //: input g0 (A) @(386,240) /sn:0 /w:[ 0 ]
  //: joint g13 (B) @(449, 246) /w:[ 2 -1 1 4 ]

endmodule

module main;    //: root_module
wire w16;    //: /sn:0 {0}(383,325)(383,335){1}
wire w13;    //: /sn:0 {0}(584,382)(594,382){1}
wire w6;    //: /sn:0 {0}(872,324)(872,334){1}
wire w7;    //: /sn:0 {0}(964,374)(954,374){1}
wire w4;    //: /sn:0 {0}(1078,378)(1088,378){1}
wire w3;    //: /sn:0 {0}(1136,446)(1136,436){1}
wire w0;    //: /sn:0 {0}(1215,373)(1205,373){1}
wire w19;    //: /sn:0 {0}(396,448)(396,438){1}
wire w18;    //: /sn:0 {0}(338,380)(348,380){1}
wire w12;    //: /sn:0 {0}(721,377)(711,377){1}
wire w10;    //: /sn:0 {0}(673,327)(673,337){1}
wire w1;    //: /sn:0 {0}(1167,323)(1167,333){1}
wire w8;    //: /sn:0 {0}(827,379)(837,379){1}
wire w17;    //: /sn:0 {0}(475,375)(465,375){1}
wire w14;    //: /sn:0 {0}(642,450)(642,440){1}
wire w11;    //: /sn:0 {0}(629,327)(629,337){1}
wire w2;    //: /sn:0 {0}(1123,323)(1123,333){1}
wire w15;    //: /sn:0 {0}(427,325)(427,335){1}
wire w5;    //: /sn:0 {0}(916,324)(916,334){1}
wire w9;    //: /sn:0 {0}(885,447)(885,437){1}
//: enddecls

  FA g3 (.A(w16), .B(w15), .Ci(w17), .Co(w18), .S(w19));   //: @(349, 336) /sz:(115, 101) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<1 Bo0<1 ]
  FA g2 (.A(w11), .B(w10), .Ci(w12), .Co(w13), .S(w14));   //: @(595, 338) /sz:(115, 101) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<1 Bo0<1 ]
  FA g1 (.A(w6), .B(w5), .Ci(w7), .Co(w8), .S(w9));   //: @(838, 335) /sz:(115, 101) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<1 Bo0<1 ]
  FA g0 (.A(w2), .B(w1), .Ci(w0), .Co(w4), .S(w3));   //: @(1089, 334) /sz:(115, 101) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<1 Bo0<1 ]

endmodule
