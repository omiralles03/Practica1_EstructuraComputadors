//: version "1.8.7"

module HA(C, S, B, A);
//: interface  /sz:(148, 128) /bd:[ Li0>A(35/128) Li1>B(102/128) Ro0<S(38/128) Ro1<C(103/128) ]
input B;    //: /sn:0 {0}(197,310)(262,310)(262,284)(288,284){1}
//: {2}(292,284)(337,284){3}
//: {4}(290,286)(290,332)(343,332){5}
input A;    //: /sn:0 {0}(198,279)(304,279){1}
//: {2}(308,279)(337,279){3}
//: {4}(306,281)(306,327)(343,327){5}
output C;    //: /sn:0 /dp:1 {0}(364,330)(448,330){1}
output S;    //: /sn:0 /dp:1 {0}(358,282)(437,282)(437,281)(447,281){1}
//: enddecls

  xor g4 (.I0(A), .I1(B), .Z(S));   //: @(348,282) /sn:0 /delay:" 6" /w:[ 3 3 0 ]
  //: output g3 (C) @(445,330) /sn:0 /w:[ 1 ]
  //: output g2 (S) @(444,281) /sn:0 /w:[ 1 ]
  //: input g1 (B) @(195,310) /sn:0 /w:[ 0 ]
  //: joint g6 (A) @(306, 279) /w:[ 2 -1 1 4 ]
  //: joint g7 (B) @(290, 284) /w:[ 2 -1 1 4 ]
  and g5 (.I0(A), .I1(B), .Z(C));   //: @(354,330) /sn:0 /delay:" 5" /w:[ 5 5 0 ]
  //: input g0 (A) @(196,279) /sn:0 /w:[ 0 ]

endmodule

module main;    //: root_module
wire w13;    //: /sn:0 {0}(823,288)(873,288)(873,287)(878,287){1}
wire w3;    //: /sn:0 /dp:1 {0}(584,215)(381,215)(381,218)(374,218){1}
wire w0;    //: /sn:0 {0}(122,184)(209,184)(209,215)(224,215){1}
wire w10;    //: /sn:0 {0}(496,277)(574,277)(574,282)(584,282){1}
wire w1;    //: /sn:0 {0}(116,282)(224,282){1}
wire w8;    //: /sn:0 {0}(734,218)(874,218)(874,224)(880,224){1}
wire w5;    //: /sn:0 {0}(374,274)(425,274)(425,376)(773,376)(773,290)(802,290){1}
wire w9;    //: /sn:0 {0}(734,283)(792,283)(792,285)(802,285){1}
//: enddecls

  led g4 (.I(w8));   //: @(887,224) /sn:0 /R:3 /w:[ 1 ] /type:0
  led g3 (.I(w13));   //: @(885,287) /sn:0 /R:3 /w:[ 1 ] /type:0
  HA g2 (.B(w1), .A(w0), .C(w5), .S(w3));   //: @(225, 180) /sz:(148, 128) /sn:0 /p:[ Li0>1 Li1>1 Ro0<0 Ro1<1 ]
  //: switch g1 (w1) @(99,282) /sn:0 /w:[ 0 ] /st:0
  //: switch g6 (w10) @(479,277) /sn:0 /w:[ 0 ] /st:0
  or g7 (.I0(w9), .I1(w5), .Z(w13));   //: @(813,288) /sn:0 /delay:" 5" /w:[ 1 1 0 ]
  HA g5 (.B(w10), .A(w3), .C(w9), .S(w8));   //: @(585, 180) /sz:(148, 128) /sn:0 /p:[ Li0>1 Li1>0 Ro0<0 Ro1<0 ]
  //: switch g0 (w0) @(105,184) /sn:0 /w:[ 0 ] /st:1

endmodule
