//: version "1.8.7"

module FA(Cout, S, Cin, B, A);
//: interface  /sz:(100, 89) /bd:[ Ti0>B(70/100) Ti1>A(27/100) Li0>Cin(31/89) Bo0<S(48/100) Ro0<Cout(32/89) ]
input B;    //: /sn:0 {0}(398,307)(450,307){1}
//: {2}(454,307)(504,307){3}
//: {4}(452,309)(452,352)(556,352){5}
input A;    //: /sn:0 {0}(556,357)(438,357)(438,284){1}
//: {2}(440,282)(490,282)(490,302)(504,302){3}
//: {4}(436,282)(398,282){5}
input Cin;    //: /sn:0 {0}(398,321)(549,321){1}
//: {2}(551,319)(551,310)(560,310){3}
//: {4}(551,323)(551,332)(556,332){5}
output Cout;    //: /sn:0 /dp:1 {0}(626,344)(659,344){1}
output S;    //: /sn:0 /dp:1 {0}(581,308)(659,308){1}
wire w14;    //: /sn:0 {0}(577,355)(596,355)(596,346)(605,346){1}
wire w11;    //: /sn:0 {0}(577,335)(596,335)(596,341)(605,341){1}
wire w2;    //: /sn:0 {0}(525,305)(537,305){1}
//: {2}(541,305)(560,305){3}
//: {4}(539,307)(539,337)(556,337){5}
//: enddecls

  and g8 (.I0(Cin), .I1(w2), .Z(w11));   //: @(567,335) /sn:0 /delay:" 3" /w:[ 5 5 0 ]
  //: output g4 (Cout) @(656,344) /sn:0 /w:[ 1 ]
  //: output g3 (S) @(656,308) /sn:0 /w:[ 1 ]
  //: input g2 (Cin) @(396,321) /sn:0 /w:[ 0 ]
  //: input g1 (B) @(396,307) /sn:0 /w:[ 0 ]
  //: joint g10 (Cin) @(551, 321) /w:[ -1 2 1 4 ]
  xor g6 (.I0(w2), .I1(Cin), .Z(S));   //: @(571,308) /sn:0 /delay:" 4" /w:[ 3 3 0 ]
  and g9 (.I0(B), .I1(A), .Z(w14));   //: @(567,355) /sn:0 /delay:" 3" /w:[ 5 0 0 ]
  or g7 (.I0(w11), .I1(w14), .Z(Cout));   //: @(616,344) /sn:0 /delay:" 3" /w:[ 1 1 0 ]
  //: joint g12 (B) @(452, 307) /w:[ 2 -1 1 4 ]
  xor g5 (.I0(A), .I1(B), .Z(w2));   //: @(515,305) /sn:0 /delay:" 4" /w:[ 3 3 0 ]
  //: joint g11 (A) @(438, 282) /w:[ 2 -1 4 1 ]
  //: input g0 (A) @(396,282) /sn:0 /w:[ 5 ]
  //: joint g13 (w2) @(539, 305) /w:[ 2 -1 1 4 ]

endmodule

module main;    //: root_module
wire [3:0] w6;    //: /sn:0 {0}(681,207)(665,207)(665,241){1}
wire w3;    //: /sn:0 {0}(560,281)(594,281){1}
wire w1;    //: /sn:0 {0}(693,283)(722,283){1}
wire [3:0] w2;    //: /sn:0 {0}(644,353)(644,326){1}
wire [3:0] w5;    //: /sn:0 {0}(608,207)(624,207)(624,241){1}
//: enddecls

  //: switch g4 (w3) @(543,281) /sn:0 /w:[ 0 ] /st:1
  led g3 (.I(w2));   //: @(644,360) /sn:0 /R:2 /w:[ 0 ] /type:2
  //: dip g2 (w6) @(719,207) /sn:0 /R:3 /w:[ 0 ] /st:3
  //: dip g1 (w5) @(570,207) /sn:0 /R:1 /w:[ 0 ] /st:11
  led g5 (.I(w1));   //: @(729,283) /sn:0 /R:3 /w:[ 1 ] /type:2
  CPA_4b g0 (.B(w6), .A(w5), .Cin(w3), .S(w2), .Cout(w1));   //: @(595, 242) /sz:(97, 83) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>1 Bo0<1 Ro0<0 ]

endmodule

module CPA_4b(S, Cin, Cout, B, A);
//: interface  /sz:(97, 83) /bd:[ Ti0>B[3:0](70/97) Ti1>A[3:0](29/97) Li0>Cin(39/83) Bo0<S[3:0](49/97) Ro0<Cout(41/83) ]
input [3:0] B;    //: /sn:0 {0}(298,170)(413,170){1}
//: {2}(414,170)(550,170){3}
//: {4}(551,170)(679,170){5}
//: {6}(680,170)(816,170){7}
//: {8}(817,170)(900,170){9}
input [3:0] A;    //: /sn:0 {0}(896,147)(774,147){1}
//: {2}(773,147)(637,147){3}
//: {4}(636,147)(508,147){5}
//: {6}(507,147)(371,147){7}
//: {8}(370,147)(299,147){9}
input Cin;    //: /sn:0 {0}(295,231)(343,231){1}
output Cout;    //: /sn:0 /dp:1 {0}(848,235)(911,235){1}
output [3:0] S;    //: /sn:0 {0}(877,326)(922,326){1}
wire w16;    //: /sn:0 {0}(658,292)(658,321)(871,321){1}
wire w13;    //: /sn:0 {0}(637,201)(637,151){1}
wire w7;    //: /sn:0 {0}(817,202)(817,174){1}
wire w4;    //: /sn:0 {0}(371,199)(371,151){1}
wire w3;    //: /sn:0 /dp:1 {0}(871,331)(529,331)(529,291){1}
wire w0;    //: /sn:0 {0}(551,200)(551,174){1}
wire w10;    //: /sn:0 {0}(680,201)(680,174){1}
wire w1;    //: /sn:0 {0}(508,200)(508,151){1}
wire w8;    //: /sn:0 /dp:1 {0}(480,232)(445,232){1}
wire w14;    //: /sn:0 /dp:1 {0}(609,233)(582,233){1}
wire w11;    //: /sn:0 /dp:1 {0}(392,290)(392,341)(871,341){1}
wire w2;    //: /sn:0 {0}(414,199)(414,174){1}
wire w15;    //: /sn:0 /dp:1 {0}(746,234)(711,234){1}
wire w5;    //: /sn:0 /dp:1 {0}(871,311)(795,311)(795,293){1}
wire w9;    //: /sn:0 {0}(774,202)(774,151){1}
//: enddecls

  FA g4 (.A(w4), .B(w2), .Cin(Cin), .S(w11), .Cout(w8));   //: @(344, 200) /sz:(100, 89) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>1 Bo0<0 Ro0<1 ]
  //: output g8 (S) @(919,326) /sn:0 /w:[ 1 ]
  //: input g3 (Cin) @(293,231) /sn:0 /w:[ 0 ]
  tran g16(.Z(w9), .I(A[3]));   //: @(774,145) /sn:0 /R:1 /w:[ 1 2 1 ] /ss:1
  tran g17(.Z(w7), .I(B[3]));   //: @(817,168) /sn:0 /R:1 /w:[ 1 7 8 ] /ss:1
  //: output g2 (Cout) @(908,235) /sn:0 /w:[ 1 ]
  //: input g1 (B) @(296,170) /sn:0 /w:[ 0 ]
  tran g10(.Z(w4), .I(A[0]));   //: @(371,145) /sn:0 /R:1 /w:[ 1 8 7 ] /ss:1
  FA g6 (.A(w13), .B(w10), .Cin(w14), .S(w16), .Cout(w15));   //: @(610, 202) /sz:(100, 89) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>0 Bo0<0 Ro0<1 ]
  FA g7 (.A(w9), .B(w7), .Cin(w15), .S(w5), .Cout(Cout));   //: @(747, 203) /sz:(100, 89) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>0 Bo0<1 Ro0<0 ]
  concat g9 (.I0(w11), .I1(w3), .I2(w16), .I3(w5), .Z(S));   //: @(876,326) /sn:0 /w:[ 1 0 1 0 0 ] /dr:0
  tran g12(.Z(w1), .I(A[1]));   //: @(508,145) /sn:0 /R:1 /w:[ 1 6 5 ] /ss:1
  FA g5 (.A(w1), .B(w0), .Cin(w8), .S(w3), .Cout(w14));   //: @(481, 201) /sz:(100, 89) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>0 Bo0<1 Ro0<1 ]
  tran g11(.Z(w2), .I(B[0]));   //: @(414,168) /sn:0 /R:1 /w:[ 1 1 2 ] /ss:1
  tran g14(.Z(w13), .I(A[2]));   //: @(637,145) /sn:0 /R:1 /w:[ 1 4 3 ] /ss:1
  //: input g0 (A) @(297,147) /sn:0 /w:[ 9 ]
  tran g15(.Z(w10), .I(B[2]));   //: @(680,168) /sn:0 /R:1 /w:[ 1 5 6 ] /ss:1
  tran g13(.Z(w0), .I(B[1]));   //: @(551,168) /sn:0 /R:1 /w:[ 1 3 4 ] /ss:1

endmodule
