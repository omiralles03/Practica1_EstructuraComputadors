//: version "1.8.7"

module HA(C, S, B, A);
//: interface  /sz:(97, 93) /bd:[ Li0>B(65/93) Li1>A(25/93) Ro0<C(66/93) Ro1<S(25/93) ]
input B;    //: /sn:0 {0}(229,171)(256,171){1}
//: {2}(260,171)(287,171){3}
//: {4}(258,173)(258,197)(287,197){5}
input A;    //: /sn:0 {0}(228,146)(243,146)(243,166)(272,166){1}
//: {2}(276,166)(287,166){3}
//: {4}(274,168)(274,192)(287,192){5}
output C;    //: /sn:0 /dp:1 {0}(308,195)(341,195){1}
output S;    //: /sn:0 /dp:1 {0}(308,169)(340,169){1}
//: enddecls

  xor g4 (.I0(A), .I1(B), .Z(S));   //: @(298,169) /sn:0 /delay:" 4" /w:[ 3 3 0 ]
  //: output g3 (C) @(338,195) /sn:0 /w:[ 1 ]
  //: output g2 (S) @(337,169) /sn:0 /w:[ 1 ]
  //: input g1 (B) @(227,171) /sn:0 /w:[ 0 ]
  //: joint g6 (A) @(274, 166) /w:[ 2 -1 1 4 ]
  //: joint g7 (B) @(258, 171) /w:[ 2 -1 1 4 ]
  and g5 (.I0(A), .I1(B), .Z(C));   //: @(298,195) /sn:0 /delay:" 3" /w:[ 5 5 0 ]
  //: input g0 (A) @(226,146) /sn:0 /w:[ 0 ]

endmodule

module SUB_16b(Cin, B, A, Cout, S);
//: interface  /sz:(104, 93) /bd:[ Ti0>A[15:0](28/104) Ti1>B[15:0](66/104) Li0>Cin(45/93) Bi0>S[15:0](51/104) Ri0>Cout(45/93) ]
input [15:0] B;    //: /sn:0 /dp:1 {0}(390,184)(390,201){1}
input [15:0] A;    //: /sn:0 {0}(351,187)(351,237){1}
input Cin;    //: /sn:0 {0}(297,285)(320,285){1}
output Cout;    //: /sn:0 {0}(451,285)(425,285){1}
output [15:0] S;    //: /sn:0 {0}(373,368)(373,331){1}
wire [15:0] w5;    //: /sn:0 /dp:1 {0}(390,217)(390,237){1}
//: enddecls

  //: input g4 (Cin) @(295,285) /sn:0 /w:[ 0 ]
  //: input g3 (B) @(390,182) /sn:0 /R:3 /w:[ 0 ]
  not g2 (.I(B), .Z(w5));   //: @(390,207) /sn:0 /R:3 /w:[ 1 0 ]
  //: input g1 (A) @(351,185) /sn:0 /R:3 /w:[ 0 ]
  //: output g6 (Cout) @(448,285) /sn:0 /w:[ 0 ]
  //: output g5 (S) @(373,365) /sn:0 /R:3 /w:[ 0 ]
  CPA_16b g0 (.A(A), .B(w5), .Cin(Cin), .S(S), .Cout(Cout));   //: @(321, 238) /sz:(103, 92) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>1 Bo0<1 Ro0<1 ]

endmodule

module CPA_16b(Cin, B, S, A, Cout);
//: interface  /sz:(103, 92) /bd:[ Ti0>B[15:0](69/103) Ti1>A[15:0](30/103) Li0>Cin(47/92) Bo0<S[15:0](52/103) Ro0<Cout(47/92) ]
input [15:0] B;    //: /sn:0 /dp:1 {0}(299,175)(411,175){1}
//: {2}(412,175)(540,175){3}
//: {4}(541,175)(666,175){5}
//: {6}(667,175)(798,175){7}
//: {8}(799,175)(905,175){9}
input [15:0] A;    //: /sn:0 {0}(907,145)(758,145){1}
//: {2}(757,145)(626,145){3}
//: {4}(625,145)(500,145){5}
//: {6}(499,145)(371,145){7}
//: {8}(370,145)(300,145){9}
input Cin;    //: /sn:0 {0}(290,244)(341,244){1}
output Cout;    //: /sn:0 /dp:1 {0}(827,248)(896,248){1}
output [15:0] S;    //: /sn:0 /dp:1 {0}(853,330)(901,330){1}
wire [3:0] w6;    //: /sn:0 {0}(667,206)(667,179){1}
wire [3:0] w13;    //: /sn:0 {0}(799,207)(799,179){1}
wire [3:0] w7;    //: /sn:0 {0}(520,290)(520,335)(847,335){1}
wire w4;    //: /sn:0 {0}(440,245)(470,245){1}
wire [3:0] w0;    //: /sn:0 {0}(412,204)(412,179){1}
wire w12;    //: /sn:0 {0}(695,247)(728,247){1}
wire [3:0] w18;    //: /sn:0 /dp:1 {0}(847,315)(778,315)(778,292){1}
wire [3:0] w10;    //: /sn:0 /dp:1 {0}(847,345)(391,345)(391,289){1}
wire [3:0] w1;    //: /sn:0 {0}(371,204)(371,149){1}
wire w8;    //: /sn:0 {0}(569,246)(596,246){1}
wire [3:0] w17;    //: /sn:0 /dp:1 {0}(847,325)(646,325)(646,291){1}
wire [3:0] w14;    //: /sn:0 {0}(758,207)(758,149){1}
wire [3:0] w2;    //: /sn:0 {0}(541,205)(541,179){1}
wire [3:0] w5;    //: /sn:0 {0}(500,205)(500,149){1}
wire [3:0] w9;    //: /sn:0 {0}(626,206)(626,149){1}
//: enddecls

  tran g4(.Z(w1), .I(A[3:0]));   //: @(371,143) /sn:0 /R:1 /w:[ 1 8 7 ] /ss:1
  tran g8(.Z(w2), .I(B[7:4]));   //: @(541,173) /sn:0 /R:1 /w:[ 1 3 4 ] /ss:1
  //: input g3 (Cin) @(288,244) /sn:0 /w:[ 0 ]
  tran g16(.Z(w14), .I(A[15:12]));   //: @(758,143) /sn:0 /R:1 /w:[ 1 2 1 ] /ss:1
  tran g17(.Z(w13), .I(B[15:12]));   //: @(799,173) /sn:0 /R:1 /w:[ 1 7 8 ] /ss:1
  CPA_4b g2 (.A(w1), .B(w0), .Cin(Cin), .S(w10), .Cout(w4));   //: @(342, 205) /sz:(97, 83) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>1 Bo0<1 Ro0<0 ]
  //: input g1 (B) @(297,175) /sn:0 /w:[ 0 ]
  CPA_4b g10 (.A(w14), .B(w13), .Cin(w12), .S(w18), .Cout(Cout));   //: @(729, 208) /sz:(97, 83) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>1 Bo0<1 Ro0<0 ]
  CPA_4b g6 (.A(w5), .B(w2), .Cin(w4), .S(w7), .Cout(w8));   //: @(471, 206) /sz:(97, 83) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>1 Bo0<0 Ro0<0 ]
  tran g7(.Z(w5), .I(A[7:4]));   //: @(500,143) /sn:0 /R:1 /w:[ 1 6 5 ] /ss:1
  CPA_4b g9 (.A(w9), .B(w6), .Cin(w8), .S(w17), .Cout(w12));   //: @(597, 207) /sz:(97, 83) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>1 Bo0<1 Ro0<0 ]
  concat g12 (.I0(w10), .I1(w7), .I2(w17), .I3(w18), .Z(S));   //: @(852,330) /sn:0 /w:[ 0 1 0 0 0 ] /dr:0
  tran g5(.Z(w0), .I(B[3:0]));   //: @(412,173) /sn:0 /R:1 /w:[ 1 1 2 ] /ss:1
  //: output g11 (S) @(898,330) /sn:0 /w:[ 1 ]
  tran g14(.Z(w9), .I(A[11:8]));   //: @(626,143) /sn:0 /R:1 /w:[ 1 4 3 ] /ss:1
  //: input g0 (A) @(298,145) /sn:0 /w:[ 9 ]
  tran g15(.Z(w6), .I(B[11:8]));   //: @(667,173) /sn:0 /R:1 /w:[ 1 5 6 ] /ss:1
  //: output g13 (Cout) @(893,248) /sn:0 /w:[ 1 ]

endmodule

module main;    //: root_module
supply1 w2;    //: /sn:0 {0}(526,288)(526,305)(575,305){1}
wire [15:0] w6;    //: /sn:0 /dp:1 {0}(675,227)(642,227)(642,259){1}
wire [15:0] w4;    //: /sn:0 /dp:1 {0}(575,228)(604,228)(604,259){1}
wire w1;    //: /sn:0 {0}(716,305)(681,305){1}
wire [15:0] w5;    //: /sn:0 {0}(627,377)(627,354){1}
//: enddecls

  //: dip g3 (w6) @(713,227) /sn:0 /R:3 /w:[ 0 ] /st:5
  //: dip g2 (w4) @(537,228) /sn:0 /R:1 /w:[ 0 ] /st:10
  led g1 (.I(w5));   //: @(627,384) /sn:0 /R:2 /w:[ 0 ] /type:3
  SUB_16b g6 (.B(w6), .A(w4), .Cin(w2), .S(w5), .Cout(w1));   //: @(576, 260) /sz:(104, 93) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>1 Bi0>1 Ri0>1 ]
  led g5 (.I(w1));   //: @(723,305) /sn:0 /R:3 /w:[ 0 ] /type:2
  //: supply1 g0 (w2) @(537,288) /sn:0 /w:[ 0 ]

endmodule

module FA(Cout, S, Cin, B, A);
//: interface  /sz:(100, 89) /bd:[ Ti0>B(70/100) Ti1>A(27/100) Li0>Cin(42/89) Bo0<S(47/100) Ro0<Cout(43/89) ]
input B;    //: /sn:0 {0}(413,322)(511,322){1}
input A;    //: /sn:0 {0}(409,282)(511,282){1}
input Cin;    //: /sn:0 {0}(407,238)(670,238){1}
output Cout;    //: /sn:0 {0}(871,287)(826,287){1}
output S;    //: /sn:0 /dp:1 {0}(769,243)(873,243){1}
wire w3;    //: /sn:0 {0}(610,323)(796,323)(796,289)(805,289){1}
wire w0;    //: /sn:0 /dp:1 {0}(805,284)(769,284){1}
wire w2;    //: /sn:0 {0}(610,282)(670,282){1}
//: enddecls

  //: output g4 (Cout) @(868,287) /sn:0 /w:[ 0 ]
  //: output g3 (S) @(870,243) /sn:0 /w:[ 1 ]
  //: input g2 (Cin) @(405,238) /sn:0 /w:[ 0 ]
  //: input g1 (B) @(411,322) /sn:0 /w:[ 0 ]
  HA g6 (.B(Cin), .A(w2), .C(w0), .S(S));   //: @(671, 218) /sz:(97, 93) /sn:0 /p:[ Li0>1 Li1>1 Ro0<1 Ro1<0 ]
  or g7 (.I0(w0), .I1(w3), .Z(Cout));   //: @(816,287) /sn:0 /delay:" 3" /w:[ 0 1 1 ]
  HA g5 (.B(B), .A(A), .C(w3), .S(w2));   //: @(512, 257) /sz:(97, 93) /sn:0 /p:[ Li0>1 Li1>1 Ro0<0 Ro1<0 ]
  //: input g0 (A) @(407,282) /sn:0 /w:[ 0 ]

endmodule

module CPA_4b(S, Cin, Cout, B, A);
//: interface  /sz:(97, 83) /bd:[ Ti0>A[3:0](29/97) Ti1>B[3:0](70/97) Li0>Cin(39/83) Bo0<S[3:0](49/97) Ro0<Cout(40/83) ]
input [3:0] B;    //: /sn:0 {0}(298,170)(413,170){1}
//: {2}(414,170)(550,170){3}
//: {4}(551,170)(679,170){5}
//: {6}(680,170)(816,170){7}
//: {8}(817,170)(900,170){9}
input [3:0] A;    //: /sn:0 {0}(896,147)(774,147){1}
//: {2}(773,147)(637,147){3}
//: {4}(636,147)(508,147){5}
//: {6}(507,147)(371,147){7}
//: {8}(370,147)(299,147){9}
input Cin;    //: /sn:0 {0}(295,231)(343,231){1}
output Cout;    //: /sn:0 /dp:1 {0}(848,235)(911,235){1}
output [3:0] S;    //: /sn:0 {0}(877,326)(922,326){1}
wire w16;    //: /sn:0 /dp:1 {0}(794,282)(794,311)(871,311){1}
wire w13;    //: /sn:0 {0}(817,191)(817,174){1}
wire w6;    //: /sn:0 {0}(680,190)(680,174){1}
wire w7;    //: /sn:0 {0}(528,280)(528,331)(871,331){1}
wire w4;    //: /sn:0 {0}(445,232)(480,232){1}
wire w3;    //: /sn:0 {0}(551,189)(551,174){1}
wire w0;    //: /sn:0 {0}(414,188)(414,174){1}
wire w12;    //: /sn:0 {0}(711,234)(746,234){1}
wire w10;    //: /sn:0 {0}(871,341)(391,341)(391,279){1}
wire w1;    //: /sn:0 {0}(371,188)(371,151){1}
wire w8;    //: /sn:0 {0}(582,233)(609,233){1}
wire w17;    //: /sn:0 {0}(871,321)(657,321)(657,281){1}
wire w14;    //: /sn:0 {0}(774,191)(774,151){1}
wire w5;    //: /sn:0 {0}(508,189)(508,151){1}
wire w9;    //: /sn:0 {0}(637,190)(637,151){1}
//: enddecls

  //: output g8 (S) @(919,326) /sn:0 /w:[ 1 ]
  FA g4 (.A(w1), .B(w0), .Cin(Cin), .S(w10), .Cout(w4));   //: @(344, 189) /sz:(100, 89) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>1 Bo0<1 Ro0<0 ]
  tran g16(.Z(w14), .I(A[3]));   //: @(774,145) /sn:0 /R:1 /w:[ 1 2 1 ] /ss:1
  //: input g3 (Cin) @(293,231) /sn:0 /w:[ 0 ]
  tran g17(.Z(w13), .I(B[3]));   //: @(817,168) /sn:0 /R:1 /w:[ 1 7 8 ] /ss:1
  //: output g2 (Cout) @(908,235) /sn:0 /w:[ 1 ]
  //: input g1 (B) @(296,170) /sn:0 /w:[ 0 ]
  tran g10(.Z(w1), .I(A[0]));   //: @(371,145) /sn:0 /R:1 /w:[ 1 8 7 ] /ss:1
  FA g6 (.A(w9), .B(w6), .Cin(w8), .S(w17), .Cout(w12));   //: @(610, 191) /sz:(100, 89) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>1 Bo0<1 Ro0<0 ]
  concat g9 (.I0(w10), .I1(w7), .I2(w17), .I3(w16), .Z(S));   //: @(876,326) /sn:0 /w:[ 0 1 0 1 0 ] /dr:0
  FA g7 (.A(w14), .B(w13), .Cin(w12), .S(w16), .Cout(Cout));   //: @(747, 192) /sz:(100, 89) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>1 Bo0<0 Ro0<0 ]
  tran g12(.Z(w5), .I(A[1]));   //: @(508,145) /sn:0 /R:1 /w:[ 1 6 5 ] /ss:1
  tran g14(.Z(w9), .I(A[2]));   //: @(637,145) /sn:0 /R:1 /w:[ 1 4 3 ] /ss:1
  tran g11(.Z(w0), .I(B[0]));   //: @(414,168) /sn:0 /R:1 /w:[ 1 1 2 ] /ss:1
  FA g5 (.A(w5), .B(w3), .Cin(w4), .S(w7), .Cout(w8));   //: @(481, 190) /sz:(100, 89) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>1 Bo0<0 Ro0<0 ]
  tran g15(.Z(w6), .I(B[2]));   //: @(680,168) /sn:0 /R:1 /w:[ 1 5 6 ] /ss:1
  //: input g0 (A) @(297,147) /sn:0 /w:[ 9 ]
  tran g13(.Z(w3), .I(B[1]));   //: @(551,168) /sn:0 /R:1 /w:[ 1 3 4 ] /ss:1

endmodule
