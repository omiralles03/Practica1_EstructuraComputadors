//: version "1.8.7"

module PFA(B, S, A, Gi, Pi, Cin);
//: interface  /sz:(223, 151) /bd:[ Ti0>A(76/223) Ti1>B(147/223) Li0>Cin(73/151) Ro0<S(36/151) Ro1<Gi(113/151) Ro2<Pi(74/151) ]
input B;    //: /sn:0 {0}(312,108)(254,108){1}
//: {2}(250,108)(207,108){3}
//: {4}(252,110)(252,153){5}
//: {6}(254,155)(405,155){7}
//: {8}(252,157)(252,183)(404,183){9}
output Gi;    //: /sn:0 {0}(425,181)(453,181){1}
input A;    //: /sn:0 {0}(207,98)(281,98){1}
//: {2}(285,98)(302,98)(302,103)(312,103){3}
//: {4}(283,100)(283,148){5}
//: {6}(285,150)(405,150){7}
//: {8}(283,152)(283,178)(404,178){9}
input Cin;    //: /sn:0 {0}(199,136)(227,136)(227,127)(403,127){1}
output Pi;    //: /sn:0 /dp:1 {0}(426,153)(453,153){1}
output S;    //: /sn:0 /dp:1 {0}(424,125)(449,125){1}
wire w2;    //: /sn:0 {0}(333,106)(400,106)(400,122)(403,122){1}
//: enddecls

  //: input g8 (B) @(205,108) /sn:0 /w:[ 3 ]
  //: joint g4 (A) @(283, 98) /w:[ 2 -1 1 4 ]
  and g3 (.I0(A), .I1(B), .Z(Gi));   //: @(415,181) /sn:0 /delay:" 5" /w:[ 9 9 0 ]
  or g2 (.I0(A), .I1(B), .Z(Pi));   //: @(416,153) /sn:0 /delay:" 5" /w:[ 7 7 0 ]
  xor g1 (.I0(w2), .I1(Cin), .Z(S));   //: @(414,125) /sn:0 /delay:" 6" /w:[ 1 1 0 ]
  //: output g10 (S) @(446,125) /sn:0 /w:[ 1 ]
  //: joint g6 (B) @(252, 108) /w:[ 1 -1 2 4 ]
  //: input g9 (A) @(205,98) /sn:0 /w:[ 0 ]
  //: joint g7 (B) @(252, 155) /w:[ 6 5 -1 8 ]
  //: output g12 (Gi) @(450,181) /sn:0 /w:[ 1 ]
  //: output g11 (Pi) @(450,153) /sn:0 /w:[ 1 ]
  //: joint g5 (A) @(283, 150) /w:[ 6 5 -1 8 ]
  xor g0 (.I0(A), .I1(B), .Z(w2));   //: @(323,106) /sn:0 /delay:" 6" /w:[ 3 0 0 ]
  //: input g13 (Cin) @(197,136) /sn:0 /w:[ 0 ]

endmodule

module main;    //: root_module
wire w6;    //: /sn:0 {0}(456,287)(502,287){1}
wire w4;    //: /sn:0 {0}(22679,3979)(22679,4000){1}
wire w0;    //: /sn:0 {0}(23023,4092)(23023,4102){1}
wire w3;    //: /sn:0 {0}(627,178)(650,178)(650,213){1}
wire w10;    //: /sn:0 /dp:1 {0}(579,213)(579,178)(548,178){1}
wire w1;    //: /sn:0 {0}(23003,4096)(23003,4106){1}
wire w14;    //: /sn:0 {0}(727,250)(752,250){1}
wire w2;    //: /sn:0 {0}(4548,148)(4538,148){1}
wire w11;    //: /sn:0 {0}(821,327)(727,327){1}
wire w5;    //: /sn:0 {0}(832,288)(727,288){1}
//: enddecls

  PFA g8 (.B(w3), .A(w10), .Cin(w6), .Pi(w5), .Gi(w11), .S(w14));   //: @(503, 214) /sz:(223, 151) /sn:0 /p:[ Ti0>1 Ti1>0 Li0>1 Ro0<1 Ro1<1 Ro2<0 ]
  //: switch g4 (w6) @(439,287) /sn:0 /w:[ 0 ] /st:1
  //: switch g3 (w2) @(4566,148) /sn:0 /R:2 /w:[ 0 ] /st:0
  //: switch g2 (w1) @(23003,4083) /sn:0 /R:3 /w:[ 0 ] /st:0
  //: switch g1 (w0) @(23023,4079) /sn:0 /R:3 /w:[ 0 ] /st:0
  led g10 (.I(w11));   //: @(828,327) /sn:0 /R:3 /w:[ 0 ] /type:3
  led g6 (.I(w14));   //: @(759,250) /sn:0 /R:3 /w:[ 1 ] /type:3
  led g7 (.I(w5));   //: @(839,288) /sn:0 /R:3 /w:[ 0 ] /type:3
  //: switch g9 (w3) @(610,178) /sn:0 /w:[ 0 ] /st:0
  //: switch g5 (w4) @(22679,3966) /sn:0 /R:3 /w:[ 0 ] /st:0
  //: switch g0 (w10) @(531,178) /sn:0 /w:[ 1 ] /st:0

endmodule
