//: version "1.8.7"

module CLL(P1, C0, G2, P2, G3, C3, P0, C4, G0, C1, G1, C2, PG, P3, GG);
//: interface  /sz:(546, 40) /bd:[ Ti0>G0(487/546) Ti1>P0(459/546) Ti2>G1(346/546) Ti3>P1(318/546) Ti4>G2(201/546) Ti5>P2(173/546) Ti6>G3(52/546) Ti7>P3(24/546) Ri0>C0(19/40) To0<C3(121/546) To1<C2(274/546) To2<C1(421/546) Lo0<C4(19/40) Bo0<GG(487/546) Bo1<PG(461/546) ]
input G2;    //: /sn:0 {0}(345,293)(345,185){1}
//: {2}(347,183)(560,183){3}
//: {4}(343,183)(269,183){5}
//: {6}(265,183)(49,183){7}
//: {8}(45,183)(-68,183){9}
//: {10}(47,185)(47,249){11}
//: {12}(267,185)(267,248){13}
output GG;    //: /sn:0 /dp:1 {0}(43,314)(43,334){1}
input C0;    //: /sn:0 /dp:9 {0}(-71,61)(170,61){1}
//: {2}(174,61)(327,61){3}
//: {4}(331,61)(442,61){5}
//: {6}(446,61)(522,61){7}
//: {8}(526,61)(560,61){9}
//: {10}(524,63)(524,246){11}
//: {12}(444,63)(444,248){13}
//: {14}(329,63)(329,248){15}
//: {16}(172,63)(172,247){17}
input P1;    //: /sn:0 {0}(162,247)(162,120){1}
//: {2}(164,118)(197,118){3}
//: {4}(201,118)(317,118){5}
//: {6}(321,118)(359,118){7}
//: {8}(363,118)(432,118){9}
//: {10}(436,118)(475,118){11}
//: {12}(479,118)(560,118){13}
//: {14}(477,120)(477,247){15}
//: {16}(434,120)(434,248){17}
//: {18}(361,120)(361,249){19}
//: {20}(319,120)(319,248){21}
//: {22}(199,120)(199,247){23}
//: {24}(160,118)(113,118){25}
//: {26}(109,118)(-19,118){27}
//: {28}(-23,118)(-69,118){29}
//: {30}(-21,120)(-21,249){31}
//: {32}(111,120)(111,249){33}
output C3;    //: /sn:0 /dp:1 {0}(348,314)(348,337){1}
output PG;    //: /sn:0 /dp:1 {0}(109,270)(109,333){1}
input G0;    //: /sn:0 /dp:1 {0}(-68,97)(-18,97){1}
//: {2}(-14,97)(202,97){3}
//: {4}(206,97)(364,97){5}
//: {6}(368,97)(480,97){7}
//: {8}(484,97)(539,97){9}
//: {10}(543,97)(560,97){11}
//: {12}(541,99)(541,293){13}
//: {14}(482,99)(482,247){15}
//: {16}(366,99)(366,249){17}
//: {18}(204,99)(204,247){19}
//: {20}(-16,99)(-16,249){21}
output C4;    //: /sn:0 /dp:1 {0}(217,317)(217,337){1}
output C2;    //: /sn:0 {0}(460,337)(460,313){1}
input P3;    //: /sn:0 {0}(-31,249)(-31,204){1}
//: {2}(-29,202)(5,202){3}
//: {4}(9,202)(40,202){5}
//: {6}(44,202)(99,202){7}
//: {8}(103,202)(150,202){9}
//: {10}(154,202)(187,202){11}
//: {12}(191,202)(230,202){13}
//: {14}(234,202)(260,202){15}
//: {16}(264,202)(560,202){17}
//: {18}(262,204)(262,248){19}
//: {20}(232,204)(232,248){21}
//: {22}(189,204)(189,247){23}
//: {24}(152,204)(152,247){25}
//: {26}(101,204)(101,249){27}
//: {28}(42,204)(42,249){29}
//: {30}(7,204)(7,249){31}
//: {32}(-33,202)(-74,202){33}
input G1;    //: /sn:0 /dp:1 {0}(-67,140)(15,140){1}
//: {2}(19,140)(240,140){3}
//: {4}(244,140)(389,140){5}
//: {6}(393,140)(458,140){7}
//: {8}(462,140)(560,140){9}
//: {10}(460,142)(460,292){11}
//: {12}(391,142)(391,248){13}
//: {14}(242,142)(242,248){15}
//: {16}(17,142)(17,249){17}
input G3;    //: /sn:0 {0}(217,296)(217,222){1}
//: {2}(219,220)(560,220){3}
//: {4}(215,220)(76,220){5}
//: {6}(72,220)(-67,220){7}
//: {8}(74,222)(74,283)(50,283)(50,293){9}
input P0;    //: /sn:0 /dp:1 {0}(-67,79)(114,79){1}
//: {2}(118,79)(165,79){3}
//: {4}(169,79)(322,79){5}
//: {6}(326,79)(437,79){7}
//: {8}(441,79)(517,79){9}
//: {10}(521,79)(560,79){11}
//: {12}(519,81)(519,246){13}
//: {14}(439,81)(439,248){15}
//: {16}(324,81)(324,248){17}
//: {18}(167,81)(167,247){19}
//: {20}(116,81)(116,249){21}
output C1;    //: /sn:0 {0}(539,336)(539,314){1}
input P2;    //: /sn:0 {0}(-26,249)(-26,163){1}
//: {2}(-24,161)(10,161){3}
//: {4}(14,161)(104,161){5}
//: {6}(108,161)(155,161){7}
//: {8}(159,161)(192,161){9}
//: {10}(196,161)(235,161){11}
//: {12}(239,161)(312,161){13}
//: {14}(316,161)(354,161){15}
//: {16}(358,161)(384,161){17}
//: {18}(388,161)(560,161){19}
//: {20}(386,163)(386,248){21}
//: {22}(356,163)(356,249){23}
//: {24}(314,163)(314,248){25}
//: {26}(237,163)(237,248){27}
//: {28}(194,163)(194,247){29}
//: {30}(157,163)(157,247){31}
//: {32}(106,163)(106,249){33}
//: {34}(12,163)(12,249){35}
//: {36}(-28,161)(-72,161){37}
wire w13;    //: /sn:0 /dp:1 {0}(350,293)(350,280)(361,280)(361,270){1}
wire w6;    //: /sn:0 {0}(12,270)(12,278)(40,278)(40,293){1}
wire w7;    //: /sn:0 {0}(212,296)(212,278)(197,278)(197,268){1}
wire w4;    //: /sn:0 {0}(322,269)(322,285)(340,285)(340,293){1}
wire w0;    //: /sn:0 /dp:1 {0}(465,292)(465,284)(480,284)(480,268){1}
wire w3;    //: /sn:0 /dp:1 {0}(222,296)(222,279)(237,279)(237,269){1}
wire w12;    //: /sn:0 /dp:1 {0}(355,293)(355,285)(389,285)(389,269){1}
wire w18;    //: /sn:0 {0}(45,270)(45,293){1}
wire w10;    //: /sn:0 {0}(439,269)(439,284)(455,284)(455,292){1}
wire w21;    //: /sn:0 {0}(-23,270)(-23,283)(35,283)(35,293){1}
wire w27;    //: /sn:0 {0}(207,296)(207,285)(162,285)(162,268){1}
wire w2;    //: /sn:0 {0}(522,267)(522,283)(536,283)(536,293){1}
wire w11;    //: /sn:0 {0}(265,269)(265,287)(227,287)(227,296){1}
//: enddecls

  //: input g4 (P1) @(562,118) /sn:0 /R:2 /w:[ 13 ]
  //: input g8 (C0) @(562,61) /sn:0 /R:2 /w:[ 9 ]
  and g44 (.I0(G0), .I1(P1), .I2(P2), .I3(P3), .Z(w7));   //: @(197,258) /sn:0 /R:3 /delay:" 3" /w:[ 19 23 29 23 1 ]
  //: joint g75 (G2) @(47, 183) /w:[ 7 -1 8 10 ]
  //: input g3 (G2) @(562,183) /sn:0 /R:2 /w:[ 3 ]
  //: joint g47 (P3) @(262, 202) /w:[ 16 -1 15 18 ]
  //: joint g16 (C0) @(172, 61) /w:[ 2 -1 1 16 ]
  //: joint g17 (G0) @(541, 97) /w:[ 10 -1 9 12 ]
  //: joint g26 (C0) @(329, 61) /w:[ 4 -1 3 14 ]
  //: input g2 (P2) @(562,161) /sn:0 /R:2 /w:[ 19 ]
  //: joint g23 (P1) @(477, 118) /w:[ 12 -1 11 14 ]
  or g30 (.I0(w12), .I1(w13), .I2(G2), .I3(w4), .Z(C3));   //: @(348,304) /sn:0 /R:3 /delay:" 3" /w:[ 0 0 0 1 0 ]
  and g74 (.I0(G0), .I1(P1), .I2(P2), .I3(P3), .Z(w21));   //: @(-23,260) /sn:0 /R:3 /delay:" 3" /w:[ 21 31 0 0 0 ]
  //: input g1 (G3) @(562,220) /sn:0 /R:2 /w:[ 3 ]
  //: joint g24 (P1) @(434, 118) /w:[ 10 -1 9 16 ]
  //: joint g39 (P0) @(324, 79) /w:[ 6 -1 5 16 ]
  //: joint g77 (P3) @(7, 202) /w:[ 4 -1 3 30 ]
  and g29 (.I0(P2), .I1(G1), .Z(w12));   //: @(389,259) /sn:0 /R:3 /delay:" 3" /w:[ 21 13 1 ]
  //: joint g60 (P3) @(152, 202) /w:[ 10 -1 9 24 ]
  //: joint g51 (P3) @(232, 202) /w:[ 14 -1 13 20 ]
  or g18 (.I0(w0), .I1(G1), .I2(w10), .Z(C2));   //: @(460,303) /sn:0 /R:3 /delay:" 3" /w:[ 0 11 1 1 ]
  or g70 (.I0(G3), .I1(w18), .I2(w6), .I3(w21), .Z(GG));   //: @(43,304) /sn:0 /R:3 /delay:" 3" /w:[ 9 1 1 1 0 ]
  //: joint g82 (P1) @(-21, 118) /w:[ 27 -1 28 30 ]
  //: output g10 (C3) @(348,334) /sn:0 /R:3 /w:[ 1 ]
  //: joint g25 (P0) @(439, 79) /w:[ 8 -1 7 14 ]
  //: joint g49 (G1) @(242, 140) /w:[ 4 -1 3 14 ]
  //: joint g72 (G3) @(74, 220) /w:[ 5 -1 6 8 ]
  //: input g6 (P0) @(562,79) /sn:0 /R:2 /w:[ 11 ]
  //: joint g50 (P2) @(237, 161) /w:[ 12 -1 11 26 ]
  //: output g9 (C4) @(217,334) /sn:0 /R:3 /w:[ 1 ]
  //: input g7 (G0) @(562,97) /sn:0 /R:2 /w:[ 11 ]
  //: joint g35 (P1) @(361, 118) /w:[ 8 -1 7 18 ]
  //: joint g58 (P1) @(162, 118) /w:[ 2 -1 24 1 ]
  //: joint g68 (P2) @(106, 161) /w:[ 6 -1 5 32 ]
  and g73 (.I0(G1), .I1(P2), .I2(P3), .Z(w6));   //: @(12,260) /sn:0 /R:3 /delay:" 3" /w:[ 17 35 31 0 ]
  //: joint g56 (C0) @(524, 61) /w:[ 8 -1 7 10 ]
  //: joint g22 (G0) @(482, 97) /w:[ 8 -1 7 14 ]
  //: joint g31 (G2) @(345, 183) /w:[ 2 -1 4 1 ]
  //: joint g59 (P2) @(157, 161) /w:[ 8 -1 7 30 ]
  and g71 (.I0(P3), .I1(G2), .Z(w18));   //: @(45,260) /sn:0 /R:3 /delay:" 3" /w:[ 29 11 0 ]
  //: joint g67 (P1) @(111, 118) /w:[ 25 -1 26 32 ]
  //: joint g83 (G0) @(-16, 97) /w:[ 2 -1 1 20 ]
  //: joint g33 (P2) @(386, 161) /w:[ 18 -1 17 20 ]
  //: joint g36 (G0) @(366, 97) /w:[ 6 -1 5 16 ]
  or g41 (.I0(w11), .I1(w3), .I2(G3), .I3(w7), .I4(w27), .Z(C4));   //: @(217,307) /sn:0 /R:3 /delay:" 3" /w:[ 1 0 0 0 0 0 ]
  and g45 (.I0(C0), .I1(P0), .I2(P1), .I3(P2), .I4(P3), .Z(w27));   //: @(162,258) /sn:0 /R:3 /delay:" 3" /w:[ 17 19 0 31 25 1 ]
  //: joint g54 (P1) @(199, 118) /w:[ 4 -1 3 22 ]
  and g42 (.I0(P3), .I1(G2), .Z(w11));   //: @(265,259) /sn:0 /R:3 /delay:" 3" /w:[ 19 13 0 ]
  //: joint g52 (P3) @(189, 202) /w:[ 12 -1 11 22 ]
  //: joint g69 (P3) @(101, 202) /w:[ 8 -1 7 26 ]
  //: joint g81 (P2) @(-26, 161) /w:[ 2 -1 36 1 ]
  //: joint g40 (C0) @(444, 61) /w:[ 6 -1 5 12 ]
  //: joint g66 (P0) @(116, 79) /w:[ 2 -1 1 20 ]
  //: output g12 (C1) @(539,333) /sn:0 /R:3 /w:[ 0 ]
  and g28 (.I0(G0), .I1(P1), .I2(P2), .Z(w13));   //: @(361,260) /sn:0 /R:3 /delay:" 3" /w:[ 17 19 23 1 ]
  //: joint g34 (P2) @(356, 161) /w:[ 16 -1 15 22 ]
  //: joint g46 (G3) @(217, 220) /w:[ 2 -1 4 1 ]
  //: joint g57 (P0) @(167, 79) /w:[ 4 -1 3 18 ]
  //: input g5 (G1) @(562,140) /sn:0 /R:2 /w:[ 9 ]
  //: output g11 (C2) @(460,334) /sn:0 /R:3 /w:[ 0 ]
  or g14 (.I0(w2), .I1(G0), .Z(C1));   //: @(539,304) /sn:0 /R:3 /delay:" 3" /w:[ 1 13 1 ]
  and g19 (.I0(P1), .I1(G0), .Z(w0));   //: @(480,258) /sn:0 /R:3 /delay:" 3" /w:[ 15 15 1 ]
  //: joint g21 (G1) @(460, 140) /w:[ 8 -1 7 10 ]
  //: output g61 (PG) @(109,330) /sn:0 /R:3 /w:[ 1 ]
  and g20 (.I0(C0), .I1(P0), .I2(P1), .Z(w10));   //: @(439,259) /sn:0 /R:3 /delay:" 3" /w:[ 13 15 17 0 ]
  //: joint g32 (G1) @(391, 140) /w:[ 6 -1 5 12 ]
  //: joint g78 (P2) @(12, 161) /w:[ 4 -1 3 34 ]
  //: joint g79 (G1) @(17, 140) /w:[ 2 -1 1 16 ]
  and g63 (.I0(P0), .I1(P1), .I2(P2), .I3(P3), .Z(PG));   //: @(109,260) /sn:0 /R:3 /delay:" 3" /w:[ 21 33 33 27 0 ]
  //: input g0 (P3) @(562,202) /sn:0 /R:2 /w:[ 17 ]
  //: joint g15 (P0) @(519, 79) /w:[ 10 -1 9 12 ]
  //: joint g38 (P1) @(319, 118) /w:[ 6 -1 5 20 ]
  and g43 (.I0(G1), .I1(P2), .I2(P3), .Z(w3));   //: @(237,259) /sn:0 /R:3 /delay:" 3" /w:[ 15 27 21 1 ]
  and g27 (.I0(C0), .I1(P0), .I2(P1), .I3(P2), .Z(w4));   //: @(322,259) /sn:0 /R:3 /delay:" 3" /w:[ 15 17 21 25 0 ]
  //: joint g48 (G2) @(267, 183) /w:[ 5 -1 6 12 ]
  //: joint g37 (P2) @(314, 161) /w:[ 14 -1 13 24 ]
  //: output g62 (GG) @(43,331) /sn:0 /R:3 /w:[ 1 ]
  //: joint g55 (G0) @(204, 97) /w:[ 4 -1 3 18 ]
  //: joint g80 (P3) @(-31, 202) /w:[ 2 -1 32 1 ]
  and g13 (.I0(P0), .I1(C0), .Z(w2));   //: @(522,257) /sn:0 /R:3 /delay:" 3" /w:[ 13 11 0 ]
  //: joint g53 (P2) @(194, 161) /w:[ 10 -1 9 28 ]
  //: joint g76 (P3) @(42, 202) /w:[ 6 -1 5 28 ]

endmodule

module PFA(Cin, B, Pi, S, A, Gi);
//: interface  /sz:(99, 88) /bd:[ Ti0>A(28/99) Ti1>B(69/99) Ri0>Cin(45/88) Bo0<S(76/99) Bo1<Gi(48/99) Bo2<Pi(20/99) ]
input B;    //: /sn:0 {0}(122,203)(136,203){1}
//: {2}(140,203)(171,203){3}
//: {4}(138,205)(138,243){5}
//: {6}(140,245)(210,245){7}
//: {8}(138,247)(138,271)(210,271){9}
output Gi;    //: /sn:0 /dp:1 {0}(231,269)(254,269){1}
input A;    //: /sn:0 {0}(121,185)(143,185){1}
//: {2}(147,185)(161,185)(161,198)(171,198){3}
//: {4}(145,187)(145,238){5}
//: {6}(147,240)(210,240){7}
//: {8}(145,242)(145,266)(210,266){9}
input Cin;    //: /sn:0 {0}(122,220)(210,220){1}
output Pi;    //: /sn:0 /dp:1 {0}(231,243)(255,243){1}
output S;    //: /sn:0 /dp:1 {0}(231,218)(255,218){1}
wire w3;    //: /sn:0 /dp:1 {0}(210,215)(201,215)(201,201)(192,201){1}
//: enddecls

  //: joint g8 (B) @(138, 203) /w:[ 2 -1 1 4 ]
  xor g4 (.I0(w3), .I1(Cin), .Z(S));   //: @(221,218) /sn:0 /delay:" 4" /w:[ 0 1 0 ]
  xor g3 (.I0(A), .I1(B), .Z(w3));   //: @(182,201) /sn:0 /delay:" 4" /w:[ 3 3 1 ]
  //: input g2 (Cin) @(120,220) /sn:0 /w:[ 0 ]
  //: input g1 (B) @(120,203) /sn:0 /w:[ 0 ]
  //: joint g10 (A) @(145, 240) /w:[ 6 5 -1 8 ]
  or g6 (.I0(A), .I1(B), .Z(Pi));   //: @(221,243) /sn:0 /delay:" 3" /w:[ 7 7 0 ]
  //: joint g9 (B) @(138, 245) /w:[ 6 5 -1 8 ]
  //: joint g7 (A) @(145, 185) /w:[ 2 -1 1 4 ]
  //: output g12 (Pi) @(252,243) /sn:0 /w:[ 1 ]
  //: output g11 (S) @(252,218) /sn:0 /w:[ 1 ]
  and g5 (.I0(A), .I1(B), .Z(Gi));   //: @(221,269) /sn:0 /delay:" 3" /w:[ 9 9 0 ]
  //: input g0 (A) @(119,185) /sn:0 /w:[ 0 ]
  //: output g13 (Gi) @(251,269) /sn:0 /w:[ 1 ]

endmodule

module main;    //: root_module
wire w7;    //: /sn:0 {0}(196,273)(225,273){1}
wire [15:0] w4;    //: /sn:0 /dp:1 {0}(218,194)(255,194)(255,223){1}
wire w3;    //: /sn:0 {0}(331,272)(363,272){1}
wire w0;    //: /sn:0 {0}(281,331)(281,318){1}
wire w1;    //: /sn:0 {0}(312,331)(312,318){1}
wire [15:0] w8;    //: /sn:0 /dp:1 {0}(299,223)(299,194)(332,194){1}
wire [15:0] w5;    //: /sn:0 /dp:1 {0}(219,347)(249,347)(249,318){1}
//: enddecls

  CLA_16b g8 (.B(w8), .A(w4), .Cin(w7), .GG(w1), .PG(w0), .S(w5), .Cout(w3));   //: @(226, 224) /sz:(104, 93) /sn:0 /p:[ Ti0>0 Ti1>1 Li0>1 Bo0<1 Bo1<1 Bo2<1 Ro0<0 ]
  //: dip g4 (w8) @(370,194) /sn:0 /R:3 /w:[ 1 ] /st:15
  //: dip g3 (w4) @(180,194) /sn:0 /R:1 /w:[ 0 ] /st:255
  led g2 (.I(w3));   //: @(370,272) /sn:0 /R:3 /w:[ 1 ] /type:2
  led g1 (.I(w5));   //: @(212,347) /sn:0 /R:1 /w:[ 0 ] /type:2
  led g6 (.I(w0));   //: @(281,338) /sn:0 /R:2 /w:[ 0 ] /type:2
  led g7 (.I(w1));   //: @(312,338) /sn:0 /R:2 /w:[ 0 ] /type:2
  //: switch g5 (w7) @(179,273) /sn:0 /w:[ 0 ] /st:1

endmodule

module CLA_4b(S, Cin, B, Cout, GG, PG, A);
//: interface  /sz:(104, 92) /bd:[ Ti0>B[3:0](71/104) Ti1>A[3:0](28/104) Ri0>Cin(46/92) Lo0<Cout(47/92) Bo0<GG(85/104) Bo1<PG(56/104) Bo2<S[3:0](20/104) ]
input [3:0] B;    //: /sn:0 {0}(658,241)(633,241){1}
//: {2}(632,241)(492,241){3}
//: {4}(491,241)(347,241){5}
//: {6}(346,241)(198,241){7}
//: {8}(197,241)(102,241){9}
output GG;    //: /sn:0 {0}(612,501)(612,474){1}
input [3:0] A;    //: /sn:0 {0}(659,207)(592,207){1}
//: {2}(591,207)(451,207){3}
//: {4}(450,207)(306,207){5}
//: {6}(305,207)(157,207){7}
//: {8}(156,207)(103,207){9}
output PG;    //: /sn:0 {0}(586,501)(586,474){1}
input Cin;    //: /sn:0 {0}(743,305)(713,305){1}
//: {2}(709,305)(664,305){3}
//: {4}(711,307)(711,452)(672,452){5}
output Cout;    //: /sn:0 {0}(86,452)(124,452){1}
output [3:0] S;    //: /sn:0 {0}(86,388)(117,388){1}
wire w6;    //: /sn:0 {0}(451,260)(451,211){1}
wire w13;    //: /sn:0 {0}(149,432)(149,349){1}
wire w4;    //: /sn:0 /dp:1 {0}(205,349)(205,373)(123,373){1}
wire w0;    //: /sn:0 {0}(198,259)(198,245){1}
wire w3;    //: /sn:0 {0}(177,349)(177,432){1}
wire w22;    //: /sn:0 {0}(612,349)(612,432){1}
wire w20;    //: /sn:0 {0}(123,403)(640,403)(640,349){1}
wire w12;    //: /sn:0 {0}(326,350)(326,432){1}
wire w18;    //: /sn:0 {0}(633,259)(633,245){1}
wire w19;    //: /sn:0 {0}(592,259)(592,211){1}
wire w23;    //: /sn:0 {0}(471,432)(471,350){1}
wire w10;    //: /sn:0 {0}(246,432)(246,305)(229,305){1}
wire w21;    //: /sn:0 {0}(584,349)(584,432){1}
wire w24;    //: /sn:0 {0}(123,393)(499,393)(499,350){1}
wire w1;    //: /sn:0 {0}(157,259)(157,211){1}
wire w8;    //: /sn:0 {0}(347,260)(347,245){1}
wire w14;    //: /sn:0 {0}(399,432)(399,306)(378,306){1}
wire w2;    //: /sn:0 {0}(298,432)(298,350){1}
wire w11;    //: /sn:0 {0}(546,432)(546,306)(523,306){1}
wire w15;    //: /sn:0 {0}(443,350)(443,432){1}
wire w5;    //: /sn:0 {0}(492,260)(492,245){1}
wire w9;    //: /sn:0 {0}(306,260)(306,211){1}
wire w26;    //: /sn:0 {0}(123,383)(354,383)(354,350){1}
//: enddecls

  tran g8(.Z(w8), .I(B[2]));   //: @(347,239) /sn:0 /R:1 /w:[ 1 6 5 ] /ss:1
  PFA g4 (.A(w9), .B(w8), .Cin(w14), .S(w26), .Gi(w12), .Pi(w2));   //: @(278, 261) /sz:(99, 88) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Bo0<1 Bo1<0 Bo2<1 ]
  PFA g3 (.A(w1), .B(w0), .Cin(w10), .S(w4), .Gi(w3), .Pi(w13));   //: @(129, 260) /sz:(99, 88) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Bo0<0 Bo1<0 Bo2<1 ]
  //: joint g16 (Cin) @(711, 305) /w:[ 1 -1 2 4 ]
  //: output g17 (S) @(89,388) /sn:0 /R:2 /w:[ 0 ]
  //: input g2 (Cin) @(745,305) /sn:0 /R:2 /w:[ 0 ]
  //: input g1 (B) @(100,241) /sn:0 /w:[ 9 ]
  concat g18 (.I0(w20), .I1(w24), .I2(w26), .I3(w4), .Z(S));   //: @(118,388) /sn:0 /R:2 /w:[ 0 0 0 1 1 ] /dr:1
  tran g10(.Z(w6), .I(A[1]));   //: @(451,205) /sn:0 /R:1 /w:[ 1 4 3 ] /ss:1
  tran g6(.Z(w0), .I(B[3]));   //: @(198,239) /sn:0 /R:1 /w:[ 1 8 7 ] /ss:1
  tran g7(.Z(w9), .I(A[2]));   //: @(306,205) /sn:0 /R:1 /w:[ 1 6 5 ] /ss:1
  PFA g9 (.A(w6), .B(w5), .Cin(w11), .S(w24), .Gi(w23), .Pi(w15));   //: @(423, 261) /sz:(99, 88) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Bo0<1 Bo1<1 Bo2<0 ]
  PFA g12 (.A(w19), .B(w18), .Cin(Cin), .S(w20), .Gi(w22), .Pi(w21));   //: @(564, 260) /sz:(99, 88) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>3 Bo0<1 Bo1<0 Bo2<0 ]
  tran g5(.Z(w1), .I(A[3]));   //: @(157,205) /sn:0 /R:1 /w:[ 1 8 7 ] /ss:1
  tran g11(.Z(w5), .I(B[1]));   //: @(492,239) /sn:0 /R:1 /w:[ 1 4 3 ] /ss:1
  tran g14(.Z(w18), .I(B[0]));   //: @(633,239) /sn:0 /R:1 /w:[ 1 2 1 ] /ss:1
  //: output g19 (Cout) @(89,452) /sn:0 /R:2 /w:[ 0 ]
  //: output g21 (GG) @(612,498) /sn:0 /R:3 /w:[ 0 ]
  //: output g20 (PG) @(586,498) /sn:0 /R:3 /w:[ 0 ]
  //: input g0 (A) @(101,207) /sn:0 /w:[ 9 ]
  CLL g15 (.G0(w22), .P0(w21), .G1(w23), .P1(w15), .G2(w12), .P2(w2), .G3(w3), .P3(w13), .C0(Cin), .C3(w10), .C2(w14), .C1(w11), .C4(Cout), .GG(GG), .PG(PG));   //: @(125, 433) /sz:(546, 40) /sn:0 /p:[ Ti0>1 Ti1>1 Ti2>0 Ti3>1 Ti4>1 Ti5>0 Ti6>1 Ti7>0 Ri0>5 To0<0 To1<0 To2<0 Lo0<1 Bo0<1 Bo1<1 ]
  tran g13(.Z(w19), .I(A[0]));   //: @(592,205) /sn:0 /R:1 /w:[ 1 2 1 ] /ss:1

endmodule

module CLA_16b(GG, B, Cin, S, PG, A, Cout);
//: interface  /sz:(104, 93) /bd:[ Ti0>A[15:0](29/104) Ti1>B[15:0](73/104) Li0>Cin(49/93) Bo0<S[15:0](23/104) Bo1<PG(55/104) Bo2<GG(86/104) Ro0<Cout(48/93) ]
input [15:0] B;    //: /sn:0 {0}(829,62)(735,62){1}
//: {2}(734,62)(568,62){3}
//: {4}(567,62)(404,62){5}
//: {6}(403,62)(231,62){7}
//: {8}(230,62)(147,62){9}
output GG;    //: /sn:0 {0}(752,376)(752,354){1}
input [15:0] A;    //: /sn:0 {0}(828,35)(692,35){1}
//: {2}(691,35)(525,35){3}
//: {4}(524,35)(361,35){5}
//: {6}(360,35)(188,35){7}
//: {8}(187,35)(144,35){9}
output PG;    //: /sn:0 /dp:1 {0}(722,376)(722,354){1}
input Cin;    //: /sn:0 {0}(784,317)(806,317)(806,153){1}
//: {2}(808,151)(826,151){3}
//: {4}(804,151)(769,151){5}
output Cout;    //: /sn:0 {0}(97,317)(128,317){1}
output [15:0] S;    //: /sn:0 {0}(100,246)(130,246){1}
wire w16;    //: /sn:0 {0}(418,198)(418,285){1}
wire [3:0] w6;    //: /sn:0 {0}(404,104)(404,66){1}
wire [3:0] w7;    //: /sn:0 {0}(361,104)(361,39){1}
wire [3:0] w25;    //: /sn:0 {0}(180,201)(180,231)(136,231){1}
wire w4;    //: /sn:0 {0}(720,198)(720,285){1}
wire w36;    //: /sn:0 {0}(290,285)(290,154)(265,154){1}
wire w3;    //: /sn:0 {0}(749,198)(749,285){1}
wire [3:0] w0;    //: /sn:0 {0}(735,104)(735,66){1}
wire [3:0] w20;    //: /sn:0 {0}(188,107)(188,39){1}
wire [3:0] w29;    //: /sn:0 /dp:1 {0}(136,251)(517,251)(517,198){1}
wire w37;    //: /sn:0 {0}(457,285)(457,151)(438,151){1}
wire [3:0] w19;    //: /sn:0 {0}(231,107)(231,66){1}
wire w12;    //: /sn:0 {0}(553,198)(553,285){1}
wire w10;    //: /sn:0 {0}(312,136)(312,152)(332,152){1}
wire w23;    //: /sn:0 {0}(245,201)(245,285){1}
wire w24;    //: /sn:0 {0}(216,201)(216,285){1}
wire [3:0] w31;    //: /sn:0 /dp:1 {0}(136,241)(353,241)(353,198){1}
wire [3:0] w1;    //: /sn:0 {0}(692,104)(692,39){1}
wire [3:0] w8;    //: /sn:0 {0}(525,104)(525,39){1}
wire w27;    //: /sn:0 {0}(143,137)(143,155)(159,155){1}
wire w17;    //: /sn:0 {0}(389,198)(389,285){1}
wire [3:0] w28;    //: /sn:0 /dp:1 {0}(136,261)(684,261)(684,198){1}
wire w11;    //: /sn:0 {0}(582,198)(582,285){1}
wire [3:0] w2;    //: /sn:0 {0}(568,104)(568,66){1}
wire w38;    //: /sn:0 {0}(624,285)(624,151)(602,151){1}
wire w26;    //: /sn:0 {0}(480,131)(480,152)(496,152){1}
wire w9;    //: /sn:0 {0}(639,131)(639,152)(663,152){1}
//: enddecls

  led g4 (.I(w9));   //: @(639,124) /sn:0 /w:[ 0 ] /type:0
  CLL g8 (.P3(w24), .G3(w23), .P2(w17), .G2(w16), .P1(w12), .G1(w11), .P0(w4), .G0(w3), .C0(Cin), .C1(w38), .C2(w37), .C3(w36), .C4(Cout), .PG(PG), .GG(GG));   //: @(129, 286) /sz:(654, 67) /sn:0 /p:[ Ti0>1 Ti1>1 Ti2>1 Ti3>1 Ti4>1 Ti5>1 Ti6>1 Ti7>1 Ri0>0 To0<0 To1<0 To2<0 Lo0<1 Bo0<1 Bo1<1 ]
  concat g16 (.I0(w28), .I1(w29), .I2(w31), .I3(w25), .Z(S));   //: @(131,246) /sn:0 /R:2 /w:[ 0 0 0 1 1 ] /dr:1
  CLA_4b g3 (.A(w8), .B(w2), .Cin(w38), .Cout(w26), .S(w29), .PG(w12), .GG(w11));   //: @(497, 105) /sz:(104, 92) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Lo0<1 Bo0<1 Bo1<0 Bo2<0 ]
  //: output g17 (GG) @(752,373) /sn:0 /R:3 /w:[ 0 ]
  CLA_4b g2 (.A(w1), .B(w0), .Cin(Cin), .Cout(w9), .S(w28), .PG(w4), .GG(w3));   //: @(664, 105) /sz:(104, 92) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>5 Lo0<1 Bo0<1 Bo1<0 Bo2<0 ]
  tran g23(.Z(w7), .I(A[11:8]));   //: @(361,33) /sn:0 /R:1 /w:[ 1 6 5 ] /ss:1
  tran g24(.Z(w20), .I(A[15:12]));   //: @(188,33) /sn:0 /R:1 /w:[ 1 8 7 ] /ss:1
  //: input g1 (B) @(831,62) /sn:0 /R:2 /w:[ 0 ]
  tran g18(.Z(w1), .I(A[3:0]));   //: @(692,33) /sn:0 /R:1 /w:[ 1 2 1 ] /ss:1
  tran g25(.Z(w19), .I(B[15:12]));   //: @(231,60) /sn:0 /R:1 /w:[ 1 8 7 ] /ss:1
  led g10 (.I(w26));   //: @(480,124) /sn:0 /w:[ 0 ] /type:0
  //: input g6 (Cin) @(828,151) /sn:0 /R:2 /w:[ 3 ]
  CLA_4b g9 (.A(w20), .B(w19), .Cin(w36), .Cout(w27), .S(w25), .PG(w24), .GG(w23));   //: @(160, 108) /sz:(104, 92) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Lo0<1 Bo0<0 Bo1<0 Bo2<0 ]
  CLA_4b g7 (.A(w7), .B(w6), .Cin(w37), .Cout(w10), .S(w31), .PG(w17), .GG(w16));   //: @(333, 105) /sz:(104, 92) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Lo0<1 Bo0<1 Bo1<0 Bo2<0 ]
  tran g22(.Z(w6), .I(B[11:8]));   //: @(404,60) /sn:0 /R:1 /w:[ 1 6 5 ] /ss:1
  led g12 (.I(w27));   //: @(143,130) /sn:0 /w:[ 0 ] /type:0
  //: output g14 (S) @(103,246) /sn:0 /R:2 /w:[ 0 ]
  led g11 (.I(w10));   //: @(312,129) /sn:0 /w:[ 0 ] /type:0
  //: joint g5 (Cin) @(806, 151) /w:[ 2 -1 4 1 ]
  tran g21(.Z(w2), .I(B[7:4]));   //: @(568,60) /sn:0 /R:1 /w:[ 1 4 3 ] /ss:1
  tran g19(.Z(w0), .I(B[3:0]));   //: @(735,60) /sn:0 /R:1 /w:[ 1 2 1 ] /ss:1
  tran g20(.Z(w8), .I(A[7:4]));   //: @(525,33) /sn:0 /R:1 /w:[ 1 4 3 ] /ss:1
  //: output g15 (PG) @(722,373) /sn:0 /R:3 /w:[ 0 ]
  //: input g0 (A) @(830,35) /sn:0 /R:2 /w:[ 0 ]
  //: output g13 (Cout) @(100,317) /sn:0 /R:2 /w:[ 0 ]

endmodule
