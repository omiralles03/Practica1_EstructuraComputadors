//: version "1.8.7"

module HA(C, S, B, A);
//: interface  /sz:(97, 93) /bd:[ Li0>B(65/93) Li1>A(25/93) Ro0<C(66/93) Ro1<S(25/93) ]
input B;    //: /sn:0 {0}(229,171)(256,171){1}
//: {2}(260,171)(287,171){3}
//: {4}(258,173)(258,197)(287,197){5}
input A;    //: /sn:0 {0}(228,146)(243,146)(243,166)(272,166){1}
//: {2}(276,166)(287,166){3}
//: {4}(274,168)(274,192)(287,192){5}
output C;    //: /sn:0 /dp:1 {0}(308,195)(341,195){1}
output S;    //: /sn:0 /dp:1 {0}(308,169)(340,169){1}
//: enddecls

  xor g4 (.I0(A), .I1(B), .Z(S));   //: @(298,169) /sn:0 /delay:" 4" /w:[ 3 3 0 ]
  //: output g3 (C) @(338,195) /sn:0 /w:[ 1 ]
  //: output g2 (S) @(337,169) /sn:0 /w:[ 1 ]
  //: input g1 (B) @(227,171) /sn:0 /w:[ 0 ]
  //: joint g6 (A) @(274, 166) /w:[ 2 -1 1 4 ]
  //: joint g7 (B) @(258, 171) /w:[ 2 -1 1 4 ]
  and g5 (.I0(A), .I1(B), .Z(C));   //: @(298,195) /sn:0 /delay:" 3" /w:[ 5 5 0 ]
  //: input g0 (A) @(226,146) /sn:0 /w:[ 0 ]

endmodule

module RCA_2b(B, S, A);
//: interface  /sz:(75, 68) /bd:[ Ti0>B[1:0](51/75) Ti1>A[1:0](23/75) Bo0<S[3:0](38/75) ]
input [1:0] B;    //: /sn:0 /dp:9 {0}(8,103)(60,103){1}
//: {2}(61,103)(124,103){3}
//: {4}(125,103)(164,103){5}
//: {6}(165,103)(219,103){7}
//: {8}(220,103)(267,103){9}
input [1:0] A;    //: /sn:0 {0}(8,79)(55,79){1}
//: {2}(56,79)(119,79){3}
//: {4}(120,79)(159,79){5}
//: {6}(160,79)(214,79){7}
//: {8}(215,79)(267,79){9}
output [3:0] S;    //: /sn:0 {0}(441,321)(412,321){1}
wire w6;    //: /sn:0 {0}(59,158)(59,336)(406,336){1}
wire w16;    //: /sn:0 {0}(335,252)(363,252)(363,306)(406,306){1}
wire w13;    //: /sn:0 {0}(215,83)(215,134){1}
wire w7;    //: /sn:0 {0}(125,107)(125,133){1}
wire w4;    //: /sn:0 {0}(56,83)(56,137){1}
wire w0;    //: /sn:0 {0}(160,83)(160,132){1}
wire w3;    //: /sn:0 /dp:1 {0}(287,280)(287,316)(406,316){1}
wire w12;    //: /sn:0 {0}(165,107)(165,132){1}
wire w18;    //: /sn:0 {0}(189,251)(223,251)(236,251){1}
wire w1;    //: /sn:0 {0}(236,211)(218,211)(218,155){1}
wire w8;    //: /sn:0 {0}(120,83)(120,133){1}
wire w17;    //: /sn:0 {0}(220,107)(220,134){1}
wire w14;    //: /sn:0 {0}(162,153)(162,183){1}
wire w2;    //: /sn:0 {0}(137,282)(137,326)(406,326){1}
wire w5;    //: /sn:0 {0}(61,107)(61,137){1}
wire w9;    //: /sn:0 {0}(122,154)(122,183){1}
//: enddecls

  tran g4(.Z(w4), .I(A[0]));   //: @(56,77) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:1
  and g8 (.I0(w7), .I1(w8), .Z(w9));   //: @(122,144) /sn:0 /R:3 /delay:" 3" /w:[ 1 1 0 ]
  and g3 (.I0(w4), .I1(w5), .Z(w6));   //: @(59,148) /sn:0 /R:3 /delay:" 3" /w:[ 1 1 0 ]
  tran g16(.Z(w13), .I(A[1]));   //: @(215,77) /sn:0 /R:1 /w:[ 0 7 8 ] /ss:1
  tran g17(.Z(w17), .I(B[1]));   //: @(220,101) /sn:0 /R:1 /w:[ 0 7 8 ] /ss:1
  HA g2 (.A(w9), .B(w14), .S(w2), .C(w18));   //: @(95, 184) /sz:(93, 97) /sn:0 /p:[ Ti0>1 Ti1>1 Bo0<0 Ro0<0 ]
  //: input g1 (B) @(6,103) /sn:0 /w:[ 0 ]
  tran g10(.Z(w0), .I(A[0]));   //: @(160,77) /sn:0 /R:1 /w:[ 0 5 6 ] /ss:1
  concat g6 (.I0(w6), .I1(w2), .I2(w3), .I3(w16), .Z(S));   //: @(411,321) /sn:0 /w:[ 1 1 1 1 1 ] /dr:0
  //: output g7 (S) @(438,321) /sn:0 /w:[ 0 ]
  and g9 (.I0(w12), .I1(w0), .Z(w14));   //: @(162,143) /sn:0 /R:3 /delay:" 3" /w:[ 1 1 0 ]
  tran g12(.Z(w8), .I(A[1]));   //: @(120,77) /sn:0 /R:1 /w:[ 0 3 4 ] /ss:1
  tran g5(.Z(w5), .I(B[0]));   //: @(61,101) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:1
  tran g11(.Z(w12), .I(B[1]));   //: @(165,101) /sn:0 /R:1 /w:[ 0 5 6 ] /ss:1
  HA g14 (.A(w18), .B(w1), .S(w3), .C(w16));   //: @(237, 186) /sz:(97, 93) /sn:0 /p:[ Li0>1 Li1>0 Bo0<0 Ro0<0 ]
  //: input g0 (A) @(6,79) /sn:0 /w:[ 0 ]
  and g15 (.I0(w13), .I1(w17), .Z(w1));   //: @(218,145) /sn:0 /R:3 /delay:" 3" /w:[ 1 1 1 ]
  tran g13(.Z(w7), .I(B[0]));   //: @(125,101) /sn:0 /R:1 /w:[ 0 3 4 ] /ss:1

endmodule

module main;    //: root_module
wire [1:0] w4;    //: /sn:0 /dp:1 {0}(111,100)(134,100)(134,121){1}
wire [3:0] w3;    //: /sn:0 {0}(149,208)(149,191){1}
wire [1:0] w2;    //: /sn:0 /dp:1 {0}(183,100)(162,100)(162,121){1}
//: enddecls

  //: dip g3 (w4) @(73,100) /sn:0 /R:1 /w:[ 0 ] /st:2
  //: dip g2 (w2) @(221,100) /sn:0 /R:3 /w:[ 0 ] /st:1
  led g1 (.I(w3));   //: @(149,215) /sn:0 /R:2 /w:[ 0 ] /type:2
  RCA_2b g0 (.B(w2), .A(w4), .S(w3));   //: @(111, 122) /sz:(75, 68) /sn:0 /p:[ Ti0>1 Ti1>1 Bo0<1 ]

endmodule
