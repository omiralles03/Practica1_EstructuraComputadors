//: version "1.8.7"

module HA(C, S, B, A);
//: interface  /sz:(148, 128) /bd:[ Li0>B(102/128) Li1>A(35/128) Ro0<C(103/128) Ro1<S(38/128) ]
input B;    //: /sn:0 {0}(197,310)(262,310)(262,284)(288,284){1}
//: {2}(292,284)(337,284){3}
//: {4}(290,286)(290,332)(343,332){5}
input A;    //: /sn:0 {0}(198,279)(304,279){1}
//: {2}(308,279)(337,279){3}
//: {4}(306,281)(306,327)(343,327){5}
output C;    //: /sn:0 /dp:1 {0}(364,330)(448,330){1}
output S;    //: /sn:0 /dp:1 {0}(358,282)(437,282)(437,281)(447,281){1}
//: enddecls

  xor g4 (.I0(A), .I1(B), .Z(S));   //: @(348,282) /sn:0 /delay:" 6" /w:[ 3 3 0 ]
  //: output g3 (C) @(445,330) /sn:0 /w:[ 1 ]
  //: output g2 (S) @(444,281) /sn:0 /w:[ 1 ]
  //: input g1 (B) @(195,310) /sn:0 /w:[ 0 ]
  //: joint g6 (A) @(306, 279) /w:[ 2 -1 1 4 ]
  //: joint g7 (B) @(290, 284) /w:[ 2 -1 1 4 ]
  and g5 (.I0(A), .I1(B), .Z(C));   //: @(354,330) /sn:0 /delay:" 5" /w:[ 5 5 0 ]
  //: input g0 (A) @(196,279) /sn:0 /w:[ 0 ]

endmodule

module CPA(A, Ci, Co, S, B);
//: interface  /sz:(190, 97) /bd:[ Ti0>B[3:0](139/190) Ti1>A[3:0](56/190) Ri0>Ci(36/97) Lo0<Co(74/97) Bo0<S[3:0](92/190) ]
input [3:0] B;    //: /sn:0 {0}(1411,147)(1411,153)(1199,153){1}
//: {2}(1198,153)(845,153){3}
//: {4}(844,153)(423,153){5}
//: {6}(422,153)(222,153)(222,156)(62,156){7}
//: {8}(61,156)(33,156){9}
input [3:0] A;    //: /sn:0 /dp:3 {0}(78,87)(98,87){1}
//: {2}(99,87)(253,87)(253,89)(442,89){3}
//: {4}(443,89)(865,89){5}
//: {6}(866,89)(1214,89){7}
//: {8}(1215,89)(1435,89){9}
output Co;    //: /sn:0 /dp:1 {0}(1540,335)(1585,335){1}
input Ci;    //: /sn:0 {0}(204,439)(225,439)(225,391)(251,391){1}
output [3:0] S;    //: /sn:0 /dp:1 {0}(1372,606)(1486,606){1}
wire w6;    //: /sn:0 {0}(193,363)(243,363)(243,364)(251,364){1}
wire w16;    //: /sn:0 {0}(878,396)(845,396)(845,157){1}
wire w7;    //: /sn:0 {0}(544,361)(594,361)(594,359)(604,359){1}
wire w4;    //: /sn:0 {0}(62,160)(62,389)(118,389){1}
wire w25;    //: /sn:0 {0}(1297,355)(1359,355)(1359,357)(1369,357){1}
wire w3;    //: /sn:0 {0}(330,359)(340,359)(340,373)(372,373){1}
wire w0;    //: /sn:0 {0}(458,359)(443,359)(443,93){1}
wire w36;    //: /sn:0 /dp:1 {0}(1519,332)(1462,332)(1462,358)(1452,358){1}
wire w20;    //: /sn:0 {0}(1366,601)(742,601)(742,395)(687,395){1}
wire w29;    //: /sn:0 {0}(1452,391)(1462,391)(1462,500)(1283,500)(1283,621)(1366,621){1}
wire w18;    //: /sn:0 {0}(965,390)(1011,390)(1011,312)(1143,312)(1143,330)(1151,330){1}
wire w12;    //: /sn:0 /dp:1 {0}(785,349)(697,349)(697,363)(687,363){1}
wire w10;    //: /sn:0 {0}(544,400)(576,400)(576,313)(761,313)(761,354)(785,354){1}
wire w23;    //: /sn:0 {0}(1223,354)(1215,354)(1215,93){1}
wire w21;    //: /sn:0 {0}(1111,393)(1146,393)(1146,611)(1366,611){1}
wire w24;    //: /sn:0 {0}(1223,392)(1199,392)(1199,157){1}
wire w1;    //: /sn:0 {0}(458,399)(423,399)(423,157){1}
wire w32;    //: /sn:0 {0}(806,352)(827,352)(827,473)(1019,473)(1019,396)(1035,396){1}
wire w8;    //: /sn:0 /dp:1 {0}(372,378)(359,378)(359,327)(204,327)(204,391)(193,391){1}
wire w17;    //: /sn:0 {0}(965,355)(1035,355){1}
wire w27;    //: /sn:0 {0}(1366,591)(372,591)(372,390)(330,390){1}
wire w35;    //: /sn:0 {0}(1172,328)(1184,328)(1184,438)(1346,438)(1346,393)(1369,393){1}
wire w2;    //: /sn:0 /dp:1 {0}(1151,325)(1121,325)(1121,359)(1111,359){1}
wire w15;    //: /sn:0 {0}(878,356)(866,356)(866,93){1}
wire w5;    //: /sn:0 {0}(99,91)(99,361)(118,361){1}
wire w9;    //: /sn:0 {0}(393,376)(403,376)(403,455)(586,455)(586,400)(604,400){1}
wire w26;    //: /sn:0 {0}(1297,393)(1325,393)(1325,299)(1500,299)(1500,337)(1519,337){1}
//: enddecls

  //: input g4 (A) @(76,87) /sn:0 /w:[ 0 ]
  HA g8 (.B(w16), .A(w15), .C(w18), .S(w17));   //: @(879, 335) /sz:(85, 77) /sn:0 /p:[ Li0>0 Li1>0 Ro0<0 Ro1<0 ]
  //: input g3 (Ci) @(202,439) /sn:0 /w:[ 0 ]
  tran g16(.Z(w4), .I(B[0]));   //: @(62,154) /sn:0 /R:1 /w:[ 0 8 7 ] /ss:1
  tran g17(.Z(w0), .I(A[1]));   //: @(443,87) /sn:0 /R:1 /w:[ 1 3 4 ] /ss:1
  or g2 (.I0(w3), .I1(w8), .Z(w9));   //: @(383,376) /sn:0 /delay:" 5" /w:[ 1 0 0 ]
  //: output g23 (Co) @(1582,335) /sn:0 /w:[ 1 ]
  HA g1 (.B(w4), .A(w5), .C(w8), .S(w6));   //: @(119, 341) /sz:(73, 70) /sn:0 /p:[ Li0>1 Li1>1 Ro0<1 Ro1<0 ]
  //: output g24 (S) @(1483,606) /sn:0 /w:[ 1 ]
  tran g18(.Z(w1), .I(B[1]));   //: @(423,151) /sn:0 /R:1 /w:[ 1 6 5 ] /ss:1
  HA g10 (.B(w24), .A(w23), .C(w26), .S(w25));   //: @(1224, 334) /sz:(72, 74) /sn:0 /p:[ Li0>0 Li1>0 Ro0<0 Ro1<0 ]
  concat g25 (.I0(w29), .I1(w21), .I2(w20), .I3(w27), .Z(S));   //: @(1371,606) /sn:0 /w:[ 1 1 0 0 0 ] /dr:0
  HA g6 (.B(w1), .A(w0), .C(w10), .S(w7));   //: @(459, 339) /sz:(84, 76) /sn:0 /p:[ Li0>0 Li1>0 Ro0<0 Ro1<0 ]
  HA g7 (.B(w9), .A(w7), .C(w12), .S(w20));   //: @(605, 338) /sz:(81, 79) /sn:0 /p:[ Li0>1 Li1>1 Ro0<1 Ro1<1 ]
  HA g9 (.B(w32), .A(w17), .C(w2), .S(w21));   //: @(1036, 334) /sz:(74, 79) /sn:0 /p:[ Li0>1 Li1>1 Ro0<1 Ro1<0 ]
  tran g22(.Z(w24), .I(B[3]));   //: @(1199,151) /sn:0 /R:1 /w:[ 1 2 1 ] /ss:1
  or g12 (.I0(w12), .I1(w10), .Z(w32));   //: @(796,352) /sn:0 /delay:" 5" /w:[ 0 1 0 ]
  //: input g5 (B) @(31,156) /sn:0 /w:[ 9 ]
  HA g11 (.B(w35), .A(w25), .C(w36), .S(w29));   //: @(1370, 339) /sz:(81, 69) /sn:0 /p:[ Li0>1 Li1>1 Ro0<1 Ro1<0 ]
  or g14 (.I0(w36), .I1(w26), .Z(Co));   //: @(1530,335) /sn:0 /delay:" 5" /w:[ 0 1 0 ]
  tran g19(.Z(w16), .I(B[2]));   //: @(845,151) /sn:0 /R:1 /w:[ 1 4 3 ] /ss:1
  tran g21(.Z(w23), .I(A[3]));   //: @(1215,87) /sn:0 /R:1 /w:[ 1 7 8 ] /ss:1
  tran g20(.Z(w15), .I(A[2]));   //: @(866,87) /sn:0 /R:1 /w:[ 1 5 6 ] /ss:1
  HA g0 (.B(Ci), .A(w6), .C(w3), .S(w27));   //: @(252, 346) /sz:(77, 61) /sn:0 /p:[ Li0>1 Li1>1 Ro0<0 Ro1<1 ]
  tran g15(.Z(w5), .I(A[0]));   //: @(99,85) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:1
  or g13 (.I0(w2), .I1(w18), .Z(w35));   //: @(1162,328) /sn:0 /delay:" 5" /w:[ 0 1 0 ]

endmodule

module main;    //: root_module
wire [3:0] w4;    //: /sn:0 {0}(795,386)(795,436)(742,436)(742,320){1}
wire w0;    //: /sn:0 {0}(553,296)(649,296){1}
wire [3:0] w3;    //: /sn:0 /dp:1 {0}(820,132)(820,167)(789,167)(789,221){1}
wire w1;    //: /sn:0 {0}(902,274)(902,258)(841,258){1}
wire [3:0] w2;    //: /sn:0 {0}(684,135)(684,179)(706,179)(706,221){1}
//: enddecls

  CPA g8 (.B(w3), .A(w2), .Ci(w1), .Co(w0), .S(w4));   //: @(650, 222) /sz:(190, 97) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<1 Bo0<1 ]
  led g4 (.I(w4));   //: @(795,379) /sn:0 /w:[ 0 ] /type:3
  //: dip g3 (w3) @(820,122) /sn:0 /w:[ 0 ] /st:7
  //: dip g2 (w2) @(684,125) /sn:0 /w:[ 0 ] /st:2
  //: switch g1 (w1) @(902,288) /sn:0 /R:1 /w:[ 0 ] /st:0
  led g0 (.I(w0));   //: @(546,296) /sn:0 /R:1 /w:[ 0 ] /type:0

endmodule
