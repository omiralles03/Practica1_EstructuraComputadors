//: version "1.8.7"

module HA(C, S, B, A);
//: interface  /sz:(97, 93) /bd:[ Li0>B(65/93) Li1>A(35/128) Ro0<C(66/93) Ro1<S(25/93) ]
input B;    //: /sn:0 {0}(229,171)(256,171){1}
//: {2}(260,171)(287,171){3}
//: {4}(258,173)(258,197)(287,197){5}
input A;    //: /sn:0 {0}(228,146)(243,146)(243,166)(272,166){1}
//: {2}(276,166)(287,166){3}
//: {4}(274,168)(274,192)(287,192){5}
output C;    //: /sn:0 /dp:1 {0}(308,195)(341,195){1}
output S;    //: /sn:0 /dp:1 {0}(308,169)(340,169){1}
//: enddecls

  xor g4 (.I0(A), .I1(B), .Z(S));   //: @(298,169) /sn:0 /delay:" 4" /w:[ 3 3 0 ]
  //: output g3 (C) @(338,195) /sn:0 /w:[ 1 ]
  //: output g2 (S) @(337,169) /sn:0 /w:[ 1 ]
  //: input g1 (B) @(227,171) /sn:0 /w:[ 0 ]
  //: joint g6 (A) @(274, 166) /w:[ 2 -1 1 4 ]
  //: joint g7 (B) @(258, 171) /w:[ 2 -1 1 4 ]
  and g5 (.I0(A), .I1(B), .Z(C));   //: @(298,195) /sn:0 /delay:" 3" /w:[ 5 5 0 ]
  //: input g0 (A) @(226,146) /sn:0 /w:[ 0 ]

endmodule

module main;    //: root_module
wire w4;    //: /sn:0 {0}(468,212)(535,212){1}
wire w0;    //: /sn:0 {0}(311,171)(369,171){1}
wire w1;    //: /sn:0 {0}(311,211)(369,211){1}
wire w5;    //: /sn:0 {0}(468,171)(535,171){1}
//: enddecls

  led g4 (.I(w5));   //: @(542,171) /sn:0 /R:3 /w:[ 1 ] /type:2
  led g3 (.I(w4));   //: @(542,212) /sn:0 /R:3 /w:[ 1 ] /type:2
  HA g2 (.A(w0), .B(w1), .S(w5), .C(w4));   //: @(370, 146) /sz:(97, 93) /sn:0 /p:[ Li0>1 Li1>1 Ro0<0 Ro1<0 ]
  //: switch g1 (w1) @(294,211) /sn:0 /w:[ 0 ] /st:0
  //: switch g0 (w0) @(294,171) /sn:0 /w:[ 0 ] /st:0

endmodule
