//: version "1.8.7"

module HA(C, S, B, A);
//: interface  /sz:(148, 128) /bd:[ Li0>A(35/128) Li1>B(102/128) Ro0<S(38/128) Ro1<C(103/128) ]
input B;    //: /sn:0 {0}(197,310)(262,310)(262,284)(288,284){1}
//: {2}(292,284)(337,284){3}
//: {4}(290,286)(290,332)(343,332){5}
input A;    //: /sn:0 {0}(198,279)(304,279){1}
//: {2}(308,279)(337,279){3}
//: {4}(306,281)(306,327)(343,327){5}
output C;    //: /sn:0 /dp:1 {0}(364,330)(448,330){1}
output S;    //: /sn:0 /dp:1 {0}(358,282)(437,282)(437,281)(447,281){1}
//: enddecls

  xor g4 (.I0(A), .I1(B), .Z(S));   //: @(348,282) /sn:0 /delay:" 6" /w:[ 3 3 0 ]
  //: output g3 (C) @(445,330) /sn:0 /w:[ 1 ]
  //: output g2 (S) @(444,281) /sn:0 /w:[ 1 ]
  //: input g1 (B) @(195,310) /sn:0 /w:[ 0 ]
  //: joint g6 (A) @(306, 279) /w:[ 2 -1 1 4 ]
  //: joint g7 (B) @(290, 284) /w:[ 2 -1 1 4 ]
  and g5 (.I0(A), .I1(B), .Z(C));   //: @(354,330) /sn:0 /delay:" 5" /w:[ 5 5 0 ]
  //: input g0 (A) @(196,279) /sn:0 /w:[ 0 ]

endmodule

module main;    //: root_module
wire w3;    //: /sn:0 /dp:1 {0}(459,278)(379,278)(379,274)(374,274){1}
wire w0;    //: /sn:0 {0}(122,184)(209,184)(209,215)(224,215){1}
wire w1;    //: /sn:0 {0}(116,282)(224,282){1}
wire w2;    //: /sn:0 {0}(374,218)(456,218)(456,220)(462,220){1}
//: enddecls

  led g4 (.I(w2));   //: @(469,220) /sn:0 /R:3 /w:[ 1 ] /type:0
  led g3 (.I(w3));   //: @(466,278) /sn:0 /R:3 /w:[ 0 ] /type:0
  HA g2 (.B(w1), .A(w0), .C(w3), .S(w2));   //: @(225, 180) /sz:(148, 128) /sn:0 /p:[ Li0>1 Li1>1 Ro0<1 Ro1<0 ]
  //: switch g1 (w1) @(99,282) /sn:0 /w:[ 0 ] /st:0
  //: switch g0 (w0) @(105,184) /sn:0 /w:[ 0 ] /st:0

endmodule
