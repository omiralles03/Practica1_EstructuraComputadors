//: version "1.8.7"

module HA(C, S, B, A);
//: interface  /sz:(148, 128) /bd:[ Li0>A(35/128) Li1>B(102/128) Ro0<S(38/128) Ro1<C(103/128) ]
input B;    //: /sn:0 {0}(197,310)(262,310)(262,284)(288,284){1}
//: {2}(292,284)(337,284){3}
//: {4}(290,286)(290,332)(343,332){5}
input A;    //: /sn:0 {0}(198,279)(304,279){1}
//: {2}(308,279)(337,279){3}
//: {4}(306,281)(306,327)(343,327){5}
output C;    //: /sn:0 /dp:1 {0}(364,330)(448,330){1}
output S;    //: /sn:0 /dp:1 {0}(358,282)(437,282)(437,281)(447,281){1}
//: enddecls

  xor g4 (.I0(A), .I1(B), .Z(S));   //: @(348,282) /sn:0 /delay:" 6" /w:[ 3 3 0 ]
  //: output g3 (C) @(445,330) /sn:0 /w:[ 1 ]
  //: output g2 (S) @(444,281) /sn:0 /w:[ 1 ]
  //: input g1 (B) @(195,310) /sn:0 /w:[ 0 ]
  //: joint g6 (A) @(306, 279) /w:[ 2 -1 1 4 ]
  //: joint g7 (B) @(290, 284) /w:[ 2 -1 1 4 ]
  and g5 (.I0(A), .I1(B), .Z(C));   //: @(354,330) /sn:0 /delay:" 5" /w:[ 5 5 0 ]
  //: input g0 (A) @(196,279) /sn:0 /w:[ 0 ]

endmodule

module RCA(S, B, A);
//: interface  /sz:(128, 112) /bd:[ Ti0>A[1:0](36/128) Ti1>B[1:0](92/128) Bo0<S(62/128) ]
input [1:0] B;    //: /sn:0 {0}(489,146)(552,146){1}
//: {2}(553,146)(610,146){3}
//: {4}(611,146)(896,146){5}
//: {6}(897,146)(961,146){7}
//: {8}(962,146)(1067,146){9}
input [1:0] A;    //: /sn:0 {0}(489,94)(547,94){1}
//: {2}(548,94)(605,94){3}
//: {4}(606,94)(891,94){5}
//: {6}(892,94)(956,94){7}
//: {8}(957,94)(1042,94){9}
output [3:0] S;    //: /sn:0 {0}(1333,501)(1283,501){1}
wire w16;    //: /sn:0 {0}(999,347)(895,347)(895,234){1}
wire w6;    //: /sn:0 {0}(606,98)(606,211){1}
wire w7;    //: /sn:0 {0}(611,150)(611,211){1}
wire w4;    //: /sn:0 {0}(553,150)(553,208){1}
wire w3;    //: /sn:0 {0}(548,98)(548,208){1}
wire w0;    //: /sn:0 {0}(892,98)(892,213){1}
wire w19;    //: /sn:0 {0}(1149,415)(1200,415)(1200,516)(1277,516){1}
wire w18;    //: /sn:0 {0}(1149,350)(1217,350)(1217,506)(1277,506){1}
wire w10;    //: /sn:0 {0}(962,150)(962,218){1}
wire w1;    //: /sn:0 {0}(897,150)(897,213){1}
wire w8;    //: /sn:0 {0}(609,232)(609,414)(662,414){1}
wire w14;    //: /sn:0 {0}(812,350)(859,350)(859,496)(1277,496){1}
wire w11;    //: /sn:0 {0}(960,239)(960,486)(1277,486){1}
wire w15;    //: /sn:0 {0}(999,414)(905,414)(905,415)(812,415){1}
wire w5;    //: /sn:0 {0}(551,229)(551,347)(662,347){1}
wire w9;    //: /sn:0 {0}(957,98)(957,218){1}
//: enddecls

  tran g8(.Z(w9), .I(A[0]));   //: @(957,92) /sn:0 /R:1 /w:[ 0 7 8 ] /ss:1
  and g4 (.I0(w6), .I1(w7), .Z(w8));   //: @(609,222) /sn:0 /R:3 /delay:" 5" /w:[ 1 1 0 ]
  concat g16 (.I0(w11), .I1(w14), .I2(w18), .I3(w19), .Z(S));   //: @(1282,501) /sn:0 /w:[ 1 1 1 1 1 ] /dr:1
  and g3 (.I0(w3), .I1(w4), .Z(w5));   //: @(551,219) /sn:0 /R:3 /delay:" 5" /w:[ 1 1 0 ]
  //: output g17 (S) @(1330,501) /sn:0 /w:[ 0 ]
  and g2 (.I0(w0), .I1(w1), .Z(w16));   //: @(895,224) /sn:0 /R:3 /delay:" 5" /w:[ 1 1 1 ]
  //: input g1 (B) @(487,146) /sn:0 /w:[ 0 ]
  tran g10(.Z(w3), .I(A[0]));   //: @(548,92) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:1
  tran g6(.Z(w0), .I(A[1]));   //: @(892,92) /sn:0 /R:1 /w:[ 0 5 6 ] /ss:1
  tran g9(.Z(w10), .I(B[0]));   //: @(962,144) /sn:0 /R:1 /w:[ 0 7 8 ] /ss:1
  tran g7(.Z(w1), .I(B[1]));   //: @(897,144) /sn:0 /R:1 /w:[ 0 5 6 ] /ss:1
  tran g12(.Z(w4), .I(B[1]));   //: @(553,144) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:1
  HA g14 (.B(w8), .A(w5), .C(w15), .S(w14));   //: @(663, 312) /sz:(148, 128) /sn:0 /p:[ Li0>1 Li1>1 Ro0<1 Ro1<0 ]
  tran g11(.Z(w6), .I(A[1]));   //: @(606,92) /sn:0 /R:1 /w:[ 0 3 4 ] /ss:1
  and g5 (.I0(w9), .I1(w10), .Z(w11));   //: @(960,229) /sn:0 /R:3 /delay:" 5" /w:[ 1 1 0 ]
  HA g15 (.B(w15), .A(w16), .C(w19), .S(w18));   //: @(1000, 312) /sz:(148, 128) /sn:0 /p:[ Li0>0 Li1>0 Ro0<0 Ro1<0 ]
  //: input g0 (A) @(487,94) /sn:0 /w:[ 0 ]
  tran g13(.Z(w7), .I(B[0]));   //: @(611,144) /sn:0 /R:1 /w:[ 0 3 4 ] /ss:1

endmodule

module main;    //: root_module
wire [3:0] w0;    //: /sn:0 {0}(409,362)(409,320){1}
wire [1:0] w3;    //: /sn:0 {0}(324,131)(324,181)(383,181)(383,206){1}
wire [1:0] w1;    //: /sn:0 /dp:1 {0}(439,206)(439,178)(496,178)(496,129){1}
//: enddecls

  led g3 (.I(w0));   //: @(409,369) /sn:0 /R:2 /w:[ 0 ] /type:3
  //: dip g2 (w1) @(496,119) /sn:0 /w:[ 1 ] /st:3
  //: dip g1 (w3) @(324,121) /sn:0 /w:[ 0 ] /st:2
  RCA g0 (.B(w1), .A(w3), .S(w0));   //: @(347, 207) /sz:(128, 112) /sn:0 /p:[ Ti0>0 Ti1>1 Bo0<1 ]

endmodule
